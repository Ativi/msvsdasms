VERSION 5.7 ;

  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ONEBITADC_0
  CLASS BLOCK ;
  FOREIGN ONEBITADC_0 ;
  ORIGIN -0.605 0.000 ;
  SIZE 14.875 BY 22.530 ;
  OBS
      LAYER pwell ;
        RECT 2.795 21.150 5.805 22.530 ;
        RECT 7.955 21.150 14.405 22.530 ;
        RECT 2.325 17.300 6.275 18.610 ;
        RECT 7.485 17.300 14.875 18.610 ;
        RECT 1.075 13.590 4.085 14.970 ;
        RECT 0.605 9.740 4.555 11.050 ;
      LAYER nwell ;
        RECT 5.160 7.560 15.480 15.120 ;
      LAYER pwell ;
        RECT 0.605 4.070 4.555 5.380 ;
        RECT 1.075 0.150 4.085 1.530 ;
      LAYER nwell ;
        RECT 5.160 0.000 13.760 7.560 ;
      LAYER li1 ;
        RECT 2.885 21.335 3.135 22.345 ;
        RECT 3.745 21.335 3.995 22.345 ;
        RECT 4.605 21.335 4.855 22.345 ;
        RECT 5.465 21.335 5.715 22.345 ;
        RECT 8.045 21.335 8.295 22.345 ;
        RECT 8.905 21.335 9.155 22.345 ;
        RECT 9.765 21.335 10.015 22.345 ;
        RECT 10.625 21.335 10.875 22.345 ;
        RECT 11.485 21.335 11.735 22.345 ;
        RECT 12.345 21.335 12.595 22.345 ;
        RECT 13.205 21.335 13.455 22.345 ;
        RECT 14.065 21.335 14.315 22.345 ;
        RECT 2.885 19.235 3.135 20.245 ;
        RECT 3.745 19.235 3.995 20.245 ;
        RECT 4.605 19.235 4.855 20.245 ;
        RECT 5.465 19.235 5.715 20.245 ;
        RECT 8.045 19.235 8.295 20.245 ;
        RECT 8.905 19.235 9.155 20.245 ;
        RECT 9.765 19.235 10.015 20.245 ;
        RECT 10.625 19.235 10.875 20.245 ;
        RECT 11.485 19.235 11.735 20.245 ;
        RECT 12.345 19.235 12.595 20.245 ;
        RECT 13.205 19.235 13.455 20.245 ;
        RECT 14.065 19.235 14.315 20.245 ;
        RECT 2.455 15.455 2.705 18.985 ;
        RECT 2.885 15.455 3.135 18.985 ;
        RECT 3.315 15.455 3.565 18.985 ;
        RECT 3.745 15.455 3.995 18.985 ;
        RECT 4.175 15.455 4.425 18.985 ;
        RECT 4.605 15.455 4.855 18.985 ;
        RECT 5.035 15.455 5.285 18.985 ;
        RECT 5.465 15.455 5.715 18.985 ;
        RECT 5.895 15.455 6.145 18.985 ;
        RECT 7.615 15.455 7.865 18.985 ;
        RECT 8.045 15.455 8.295 18.985 ;
        RECT 8.475 15.455 8.725 18.985 ;
        RECT 8.905 15.455 9.155 18.985 ;
        RECT 9.335 15.455 9.585 18.985 ;
        RECT 9.765 15.455 10.015 18.985 ;
        RECT 10.195 15.455 10.445 18.985 ;
        RECT 10.625 15.455 10.875 18.985 ;
        RECT 11.055 15.455 11.305 18.985 ;
        RECT 11.485 15.455 11.735 18.985 ;
        RECT 11.915 15.455 12.165 18.985 ;
        RECT 12.345 15.455 12.595 18.985 ;
        RECT 12.775 15.455 13.025 18.985 ;
        RECT 13.205 15.455 13.455 18.985 ;
        RECT 13.635 15.455 13.885 18.985 ;
        RECT 14.065 15.455 14.315 18.985 ;
        RECT 14.495 15.455 14.745 18.985 ;
        RECT 1.165 13.775 1.415 14.785 ;
        RECT 2.025 13.775 2.275 14.785 ;
        RECT 2.885 13.775 3.135 14.785 ;
        RECT 3.745 13.775 3.995 14.785 ;
        RECT 1.165 11.675 1.415 12.685 ;
        RECT 2.025 11.675 2.275 12.685 ;
        RECT 2.885 11.675 3.135 12.685 ;
        RECT 3.745 11.675 3.995 12.685 ;
        RECT 0.735 7.895 0.985 11.425 ;
        RECT 1.165 7.895 1.415 11.425 ;
        RECT 1.595 7.895 1.845 11.425 ;
        RECT 2.025 7.895 2.275 11.425 ;
        RECT 2.455 7.895 2.705 11.425 ;
        RECT 2.885 7.895 3.135 11.425 ;
        RECT 3.315 7.895 3.565 11.425 ;
        RECT 3.745 7.895 3.995 11.425 ;
        RECT 4.175 7.895 4.425 11.425 ;
        RECT 5.895 11.255 6.145 14.785 ;
        RECT 6.325 11.255 6.575 14.785 ;
        RECT 6.755 11.255 7.005 14.785 ;
        RECT 7.185 11.255 7.435 14.785 ;
        RECT 7.615 11.255 7.865 14.785 ;
        RECT 8.045 11.255 8.295 14.785 ;
        RECT 8.475 11.255 8.725 14.785 ;
        RECT 8.905 11.255 9.155 14.785 ;
        RECT 9.335 11.255 9.585 14.785 ;
        RECT 11.055 11.255 11.305 14.785 ;
        RECT 11.485 11.255 11.735 14.785 ;
        RECT 11.915 11.255 12.165 14.785 ;
        RECT 12.345 11.255 12.595 14.785 ;
        RECT 12.775 11.255 13.025 14.785 ;
        RECT 13.205 11.255 13.455 14.785 ;
        RECT 13.635 11.255 13.885 14.785 ;
        RECT 14.065 11.255 14.315 14.785 ;
        RECT 14.495 11.255 14.745 14.785 ;
        RECT 6.325 9.995 6.575 11.005 ;
        RECT 7.185 9.995 7.435 11.005 ;
        RECT 8.045 9.995 8.295 11.005 ;
        RECT 8.905 9.995 9.155 11.005 ;
        RECT 11.485 9.995 11.735 11.005 ;
        RECT 12.345 9.995 12.595 11.005 ;
        RECT 13.205 9.995 13.455 11.005 ;
        RECT 14.065 9.995 14.315 11.005 ;
        RECT 6.325 7.895 6.575 8.905 ;
        RECT 7.185 7.895 7.435 8.905 ;
        RECT 8.045 7.895 8.295 8.905 ;
        RECT 8.905 7.895 9.155 8.905 ;
        RECT 11.485 7.895 11.735 8.905 ;
        RECT 12.345 7.895 12.595 8.905 ;
        RECT 13.205 7.895 13.455 8.905 ;
        RECT 14.065 7.895 14.315 8.905 ;
        RECT 0.735 3.695 0.985 7.225 ;
        RECT 1.165 3.695 1.415 7.225 ;
        RECT 1.595 3.695 1.845 7.225 ;
        RECT 2.025 3.695 2.275 7.225 ;
        RECT 2.455 3.695 2.705 7.225 ;
        RECT 2.885 3.695 3.135 7.225 ;
        RECT 3.315 3.695 3.565 7.225 ;
        RECT 3.745 3.695 3.995 7.225 ;
        RECT 4.175 3.695 4.425 7.225 ;
        RECT 5.895 3.695 6.145 7.225 ;
        RECT 6.325 3.695 6.575 7.225 ;
        RECT 6.755 3.695 7.005 7.225 ;
        RECT 7.185 3.695 7.435 7.225 ;
        RECT 7.615 3.695 7.865 7.225 ;
        RECT 8.045 3.695 8.295 7.225 ;
        RECT 8.475 3.695 8.725 7.225 ;
        RECT 8.905 3.695 9.155 7.225 ;
        RECT 9.335 3.695 9.585 7.225 ;
        RECT 9.765 3.695 10.015 7.225 ;
        RECT 10.195 3.695 10.445 7.225 ;
        RECT 10.625 3.695 10.875 7.225 ;
        RECT 11.055 3.695 11.305 7.225 ;
        RECT 11.485 3.695 11.735 7.225 ;
        RECT 11.915 3.695 12.165 7.225 ;
        RECT 12.345 3.695 12.595 7.225 ;
        RECT 12.775 3.695 13.025 7.225 ;
        RECT 1.165 2.435 1.415 3.445 ;
        RECT 2.025 2.435 2.275 3.445 ;
        RECT 2.885 2.435 3.135 3.445 ;
        RECT 3.745 2.435 3.995 3.445 ;
        RECT 6.325 2.435 6.575 3.445 ;
        RECT 7.185 2.435 7.435 3.445 ;
        RECT 8.045 2.435 8.295 3.445 ;
        RECT 8.905 2.435 9.155 3.445 ;
        RECT 9.765 2.435 10.015 3.445 ;
        RECT 10.625 2.435 10.875 3.445 ;
        RECT 11.485 2.435 11.735 3.445 ;
        RECT 12.345 2.435 12.595 3.445 ;
        RECT 1.165 0.335 1.415 1.345 ;
        RECT 2.025 0.335 2.275 1.345 ;
        RECT 2.885 0.335 3.135 1.345 ;
        RECT 3.745 0.335 3.995 1.345 ;
        RECT 6.325 0.335 6.575 1.345 ;
        RECT 7.185 0.335 7.435 1.345 ;
        RECT 8.045 0.335 8.295 1.345 ;
        RECT 8.905 0.335 9.155 1.345 ;
        RECT 9.765 0.335 10.015 1.345 ;
        RECT 10.625 0.335 10.875 1.345 ;
        RECT 11.485 0.335 11.735 1.345 ;
        RECT 12.345 0.335 12.595 1.345 ;
      LAYER mcon ;
        RECT 2.925 21.755 3.095 21.925 ;
        RECT 3.785 21.755 3.955 21.925 ;
        RECT 4.645 21.755 4.815 21.925 ;
        RECT 5.505 21.755 5.675 21.925 ;
        RECT 8.085 21.755 8.255 21.925 ;
        RECT 8.945 21.755 9.115 21.925 ;
        RECT 9.805 21.755 9.975 21.925 ;
        RECT 10.665 21.755 10.835 21.925 ;
        RECT 11.525 21.755 11.695 21.925 ;
        RECT 12.385 21.755 12.555 21.925 ;
        RECT 13.245 21.755 13.415 21.925 ;
        RECT 14.105 21.755 14.275 21.925 ;
        RECT 2.925 19.655 3.095 19.825 ;
        RECT 3.785 19.655 3.955 19.825 ;
        RECT 4.645 19.655 4.815 19.825 ;
        RECT 5.505 19.655 5.675 19.825 ;
        RECT 8.085 19.655 8.255 19.825 ;
        RECT 8.945 19.655 9.115 19.825 ;
        RECT 9.805 19.655 9.975 19.825 ;
        RECT 10.665 19.655 10.835 19.825 ;
        RECT 11.525 19.655 11.695 19.825 ;
        RECT 12.385 19.655 12.555 19.825 ;
        RECT 13.245 19.655 13.415 19.825 ;
        RECT 14.105 19.655 14.275 19.825 ;
        RECT 2.495 15.875 2.665 16.045 ;
        RECT 2.925 15.455 3.095 15.625 ;
        RECT 3.355 15.875 3.525 16.045 ;
        RECT 3.785 15.455 3.955 15.625 ;
        RECT 4.215 15.875 4.385 16.045 ;
        RECT 4.645 15.455 4.815 15.625 ;
        RECT 5.075 15.875 5.245 16.045 ;
        RECT 5.505 15.455 5.675 15.625 ;
        RECT 5.935 15.875 6.105 16.045 ;
        RECT 7.655 16.295 7.825 16.465 ;
        RECT 8.085 15.455 8.255 15.625 ;
        RECT 8.515 16.295 8.685 16.465 ;
        RECT 8.945 15.875 9.115 16.045 ;
        RECT 9.375 16.295 9.545 16.465 ;
        RECT 9.805 15.875 9.975 16.045 ;
        RECT 10.235 16.295 10.405 16.465 ;
        RECT 10.665 15.455 10.835 15.625 ;
        RECT 11.095 16.295 11.265 16.465 ;
        RECT 11.525 15.455 11.695 15.625 ;
        RECT 11.955 16.295 12.125 16.465 ;
        RECT 12.385 15.875 12.555 16.045 ;
        RECT 12.815 16.295 12.985 16.465 ;
        RECT 13.245 15.875 13.415 16.045 ;
        RECT 13.675 16.295 13.845 16.465 ;
        RECT 14.105 15.455 14.275 15.625 ;
        RECT 14.535 16.295 14.705 16.465 ;
        RECT 1.205 14.195 1.375 14.365 ;
        RECT 2.065 14.195 2.235 14.365 ;
        RECT 2.925 14.195 3.095 14.365 ;
        RECT 3.785 14.195 3.955 14.365 ;
        RECT 5.935 14.195 6.105 14.365 ;
        RECT 1.205 12.095 1.375 12.265 ;
        RECT 2.065 12.095 2.235 12.265 ;
        RECT 2.925 12.095 3.095 12.265 ;
        RECT 3.785 12.095 3.955 12.265 ;
        RECT 0.775 8.315 0.945 8.485 ;
        RECT 1.205 7.895 1.375 8.065 ;
        RECT 1.635 8.315 1.805 8.485 ;
        RECT 2.065 7.895 2.235 8.065 ;
        RECT 2.495 8.315 2.665 8.485 ;
        RECT 2.925 7.895 3.095 8.065 ;
        RECT 3.355 8.315 3.525 8.485 ;
        RECT 3.785 7.895 3.955 8.065 ;
        RECT 6.365 14.615 6.535 14.785 ;
        RECT 6.795 14.195 6.965 14.365 ;
        RECT 7.225 14.615 7.395 14.785 ;
        RECT 7.655 14.195 7.825 14.365 ;
        RECT 8.085 14.615 8.255 14.785 ;
        RECT 8.515 14.195 8.685 14.365 ;
        RECT 8.945 14.615 9.115 14.785 ;
        RECT 9.375 14.195 9.545 14.365 ;
        RECT 11.095 14.195 11.265 14.365 ;
        RECT 11.525 14.615 11.695 14.785 ;
        RECT 11.955 14.195 12.125 14.365 ;
        RECT 12.385 14.615 12.555 14.785 ;
        RECT 12.815 14.195 12.985 14.365 ;
        RECT 13.245 14.615 13.415 14.785 ;
        RECT 13.675 14.195 13.845 14.365 ;
        RECT 14.105 14.615 14.275 14.785 ;
        RECT 14.535 14.195 14.705 14.365 ;
        RECT 6.365 10.415 6.535 10.585 ;
        RECT 7.225 10.415 7.395 10.585 ;
        RECT 8.085 10.415 8.255 10.585 ;
        RECT 8.945 10.415 9.115 10.585 ;
        RECT 11.525 10.415 11.695 10.585 ;
        RECT 12.385 10.415 12.555 10.585 ;
        RECT 13.245 10.415 13.415 10.585 ;
        RECT 14.105 10.415 14.275 10.585 ;
        RECT 4.215 8.315 4.385 8.485 ;
        RECT 6.365 8.315 6.535 8.485 ;
        RECT 7.225 8.315 7.395 8.485 ;
        RECT 8.085 8.315 8.255 8.485 ;
        RECT 8.945 8.315 9.115 8.485 ;
        RECT 11.525 8.315 11.695 8.485 ;
        RECT 12.385 8.315 12.555 8.485 ;
        RECT 13.245 8.315 13.415 8.485 ;
        RECT 14.105 8.315 14.275 8.485 ;
        RECT 0.775 6.635 0.945 6.805 ;
        RECT 1.205 7.055 1.375 7.225 ;
        RECT 1.635 6.635 1.805 6.805 ;
        RECT 2.065 7.055 2.235 7.225 ;
        RECT 2.495 6.635 2.665 6.805 ;
        RECT 2.925 7.055 3.095 7.225 ;
        RECT 3.355 6.635 3.525 6.805 ;
        RECT 3.785 7.055 3.955 7.225 ;
        RECT 4.215 6.635 4.385 6.805 ;
        RECT 5.935 6.215 6.105 6.385 ;
        RECT 6.365 7.055 6.535 7.225 ;
        RECT 6.795 6.215 6.965 6.385 ;
        RECT 7.225 6.635 7.395 6.805 ;
        RECT 7.655 6.215 7.825 6.385 ;
        RECT 8.085 6.635 8.255 6.805 ;
        RECT 8.515 6.215 8.685 6.385 ;
        RECT 8.945 7.055 9.115 7.225 ;
        RECT 9.375 6.215 9.545 6.385 ;
        RECT 9.805 7.055 9.975 7.225 ;
        RECT 10.235 6.215 10.405 6.385 ;
        RECT 10.665 6.635 10.835 6.805 ;
        RECT 11.095 6.215 11.265 6.385 ;
        RECT 11.525 6.635 11.695 6.805 ;
        RECT 11.955 6.215 12.125 6.385 ;
        RECT 12.385 7.055 12.555 7.225 ;
        RECT 12.815 6.215 12.985 6.385 ;
        RECT 1.205 2.855 1.375 3.025 ;
        RECT 2.065 2.855 2.235 3.025 ;
        RECT 2.925 2.855 3.095 3.025 ;
        RECT 3.785 2.855 3.955 3.025 ;
        RECT 6.365 2.855 6.535 3.025 ;
        RECT 7.225 2.855 7.395 3.025 ;
        RECT 8.085 2.855 8.255 3.025 ;
        RECT 8.945 2.855 9.115 3.025 ;
        RECT 9.805 2.855 9.975 3.025 ;
        RECT 10.665 2.855 10.835 3.025 ;
        RECT 11.525 2.855 11.695 3.025 ;
        RECT 12.385 2.855 12.555 3.025 ;
        RECT 1.205 0.755 1.375 0.925 ;
        RECT 2.065 0.755 2.235 0.925 ;
        RECT 2.925 0.755 3.095 0.925 ;
        RECT 3.785 0.755 3.955 0.925 ;
        RECT 6.365 0.755 6.535 0.925 ;
        RECT 7.225 0.755 7.395 0.925 ;
        RECT 8.085 0.755 8.255 0.925 ;
        RECT 8.945 0.755 9.115 0.925 ;
        RECT 9.805 0.755 9.975 0.925 ;
        RECT 10.665 0.755 10.835 0.925 ;
        RECT 11.525 0.755 11.695 0.925 ;
        RECT 12.385 0.755 12.555 0.925 ;
      LAYER met1 ;
        RECT 2.840 21.700 5.760 21.980 ;
        RECT 8.000 21.700 14.360 21.980 ;
        RECT 2.840 19.600 7.470 19.880 ;
        RECT 8.000 19.600 14.360 19.880 ;
        RECT 7.150 19.180 10.910 19.460 ;
        RECT 4.570 18.760 11.770 19.040 ;
        RECT 7.570 16.240 14.790 16.520 ;
        RECT 2.410 15.820 6.190 16.100 ;
        RECT 8.860 15.820 13.500 16.100 ;
        RECT 2.840 15.400 5.760 15.680 ;
        RECT 8.000 15.400 14.360 15.680 ;
        RECT 7.580 14.980 10.910 15.260 ;
        RECT 6.280 14.560 9.200 14.840 ;
        RECT 11.440 14.560 14.360 14.840 ;
        RECT 1.120 14.140 4.040 14.420 ;
        RECT 5.850 14.140 9.630 14.420 ;
        RECT 11.010 14.140 14.790 14.420 ;
        RECT 1.120 12.040 4.040 12.320 ;
        RECT 6.280 10.360 9.200 10.640 ;
        RECT 11.440 10.360 14.360 10.640 ;
        RECT 0.690 8.260 4.470 8.540 ;
        RECT 6.280 8.260 9.200 8.540 ;
        RECT 11.440 8.260 14.360 8.540 ;
        RECT 1.120 7.840 7.470 8.120 ;
        RECT 8.010 7.840 12.630 8.120 ;
        RECT 1.120 7.000 5.750 7.280 ;
        RECT 6.280 7.000 12.640 7.280 ;
        RECT 0.690 6.580 4.470 6.860 ;
        RECT 7.140 6.580 11.780 6.860 ;
        RECT 5.850 6.160 13.070 6.440 ;
        RECT 1.120 2.800 4.040 3.080 ;
        RECT 6.280 2.800 12.640 3.080 ;
        RECT 1.120 0.700 4.040 0.980 ;
        RECT 6.280 0.700 12.640 0.980 ;
      LAYER via ;
        RECT 4.600 21.710 4.860 21.970 ;
        RECT 11.480 21.710 11.740 21.970 ;
        RECT 7.180 19.610 7.440 19.870 ;
        RECT 10.620 19.610 10.880 19.870 ;
        RECT 7.180 19.190 7.440 19.450 ;
        RECT 10.620 19.190 10.880 19.450 ;
        RECT 4.600 18.770 4.860 19.030 ;
        RECT 11.480 18.770 11.740 19.030 ;
        RECT 11.480 16.250 11.740 16.510 ;
        RECT 4.600 15.830 4.860 16.090 ;
        RECT 11.910 15.830 12.170 16.090 ;
        RECT 2.880 15.410 3.140 15.670 ;
        RECT 10.620 15.410 10.880 15.670 ;
        RECT 7.610 14.990 7.870 15.250 ;
        RECT 10.620 14.990 10.880 15.250 ;
        RECT 7.610 14.570 7.870 14.830 ;
        RECT 11.910 14.570 12.170 14.830 ;
        RECT 2.880 14.150 3.140 14.410 ;
        RECT 8.040 14.150 8.300 14.410 ;
        RECT 12.340 14.150 12.600 14.410 ;
        RECT 7.610 10.370 7.870 10.630 ;
        RECT 11.480 10.370 11.740 10.630 ;
        RECT 2.880 8.270 3.140 8.530 ;
        RECT 8.040 8.270 8.300 8.530 ;
        RECT 12.340 8.270 12.600 8.530 ;
        RECT 7.180 7.850 7.440 8.110 ;
        RECT 8.040 7.850 8.300 8.110 ;
        RECT 9.760 7.850 10.020 8.110 ;
        RECT 12.340 7.850 12.600 8.110 ;
        RECT 5.460 7.010 5.720 7.270 ;
        RECT 8.900 7.010 9.160 7.270 ;
        RECT 2.880 6.590 3.140 6.850 ;
        RECT 7.180 6.590 7.440 6.850 ;
        RECT 11.480 6.590 11.740 6.850 ;
        RECT 9.760 6.170 10.020 6.430 ;
        RECT 8.900 2.810 9.160 3.070 ;
        RECT 2.880 0.710 3.140 0.970 ;
        RECT 9.760 0.710 10.020 0.970 ;
      LAYER met2 ;
        RECT 4.590 15.800 4.870 22.000 ;
        RECT 7.170 19.160 7.450 19.900 ;
        RECT 2.870 0.680 3.150 15.700 ;
        RECT 7.600 10.340 7.880 15.280 ;
        RECT 10.610 14.960 10.890 19.900 ;
        RECT 11.470 16.220 11.750 22.000 ;
        RECT 11.900 14.540 12.180 16.120 ;
        RECT 5.450 6.115 5.730 7.300 ;
        RECT 7.170 6.560 7.450 8.140 ;
        RECT 8.030 7.820 8.310 14.440 ;
        RECT 8.890 2.780 9.170 7.300 ;
        RECT 9.750 0.680 10.030 8.140 ;
        RECT 11.470 6.560 11.750 10.660 ;
        RECT 12.330 7.820 12.610 14.440 ;
      LAYER via2 ;
        RECT 5.450 6.160 5.730 6.440 ;
        RECT 8.890 6.160 9.170 6.440 ;
      LAYER met3 ;
        RECT 5.425 5.900 9.195 6.700 ;
  END
END ONEBITADC_0
END LIBRARY

