module RINGOSC_0(
    output Vin
;

endmodule 
