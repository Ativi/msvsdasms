MACRO RINGOSC
  ORIGIN 0 0 ;
  FOREIGN RINGOSC 0 0 ;
  SIZE 12.04 BY 30.24 ;
  PIN GND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 3.3 8.24 3.58 14.44 ;
      LAYER M3 ;
        RECT 8.46 8.24 8.74 14.44 ;
      LAYER M3 ;
        RECT 3.3 11.155 3.58 11.525 ;
      LAYER M2 ;
        RECT 3.44 11.2 8.6 11.48 ;
      LAYER M3 ;
        RECT 8.46 11.155 8.74 11.525 ;
      LAYER M3 ;
        RECT 5.45 23.36 5.73 29.56 ;
      LAYER M3 ;
        RECT 3.3 14.28 3.58 22.68 ;
      LAYER M2 ;
        RECT 3.44 22.54 5.59 22.82 ;
      LAYER M3 ;
        RECT 5.45 22.68 5.73 23.52 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 3.3 0.68 3.58 6.88 ;
      LAYER M3 ;
        RECT 8.46 0.68 8.74 6.88 ;
      LAYER M3 ;
        RECT 3.3 3.595 3.58 3.965 ;
      LAYER M2 ;
        RECT 3.44 3.64 8.6 3.92 ;
      LAYER M3 ;
        RECT 8.46 3.595 8.74 3.965 ;
      LAYER M3 ;
        RECT 5.45 15.8 5.73 22 ;
      LAYER M3 ;
        RECT 8.46 6.72 8.74 7.56 ;
      LAYER M2 ;
        RECT 8.17 7.42 8.6 7.7 ;
      LAYER M3 ;
        RECT 8.03 7.56 8.31 21.42 ;
      LAYER M2 ;
        RECT 5.59 21.28 8.17 21.56 ;
      LAYER M3 ;
        RECT 5.45 21.235 5.73 21.605 ;
    END
  END VDD
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 7.14 2.8 10.92 3.08 ;
      LAYER M2 ;
        RECT 7.14 12.04 10.92 12.32 ;
      LAYER M2 ;
        RECT 8.87 2.8 9.19 3.08 ;
      LAYER M3 ;
        RECT 8.89 2.94 9.17 12.18 ;
      LAYER M2 ;
        RECT 8.87 12.04 9.19 12.32 ;
      LAYER M2 ;
        RECT 4.13 22.12 7.91 22.4 ;
      LAYER M2 ;
        RECT 4.13 22.96 7.91 23.24 ;
      LAYER M2 ;
        RECT 5.86 22.12 6.18 22.4 ;
      LAYER M3 ;
        RECT 5.88 22.26 6.16 23.1 ;
      LAYER M2 ;
        RECT 5.86 22.96 6.18 23.24 ;
      LAYER M2 ;
        RECT 7.15 12.04 7.47 12.32 ;
      LAYER M3 ;
        RECT 7.17 12.18 7.45 22.26 ;
      LAYER M2 ;
        RECT 7.15 22.12 7.47 22.4 ;
    END
  END Y
  OBS 
  LAYER M2 ;
        RECT 1.12 7 4.9 7.28 ;
  LAYER M2 ;
        RECT 1.12 7.84 4.9 8.12 ;
  LAYER M2 ;
        RECT 2.85 7 3.17 7.28 ;
  LAYER M3 ;
        RECT 2.87 7.14 3.15 7.98 ;
  LAYER M2 ;
        RECT 2.85 7.84 3.17 8.12 ;
  LAYER M2 ;
        RECT 4.13 17.92 7.91 18.2 ;
  LAYER M2 ;
        RECT 4.13 27.16 7.91 27.44 ;
  LAYER M2 ;
        RECT 6.29 17.92 6.61 18.2 ;
  LAYER M3 ;
        RECT 6.31 18.06 6.59 27.3 ;
  LAYER M2 ;
        RECT 6.29 27.16 6.61 27.44 ;
  LAYER M2 ;
        RECT 4.14 7.84 4.46 8.12 ;
  LAYER M3 ;
        RECT 4.16 7.98 4.44 18.06 ;
  LAYER M2 ;
        RECT 4.14 17.92 4.46 18.2 ;
  LAYER M2 ;
        RECT 4.14 7.84 4.46 8.12 ;
  LAYER M3 ;
        RECT 4.16 7.82 4.44 8.14 ;
  LAYER M2 ;
        RECT 4.14 17.92 4.46 18.2 ;
  LAYER M3 ;
        RECT 4.16 17.9 4.44 18.22 ;
  LAYER M2 ;
        RECT 4.14 7.84 4.46 8.12 ;
  LAYER M3 ;
        RECT 4.16 7.82 4.44 8.14 ;
  LAYER M2 ;
        RECT 4.14 17.92 4.46 18.2 ;
  LAYER M3 ;
        RECT 4.16 17.9 4.44 18.22 ;
  LAYER M2 ;
        RECT 1.12 2.8 4.9 3.08 ;
  LAYER M2 ;
        RECT 1.12 12.04 4.9 12.32 ;
  LAYER M2 ;
        RECT 7.14 7 10.92 7.28 ;
  LAYER M2 ;
        RECT 7.14 7.84 10.92 8.12 ;
  LAYER M2 ;
        RECT 4.57 2.8 4.89 3.08 ;
  LAYER M3 ;
        RECT 4.59 2.94 4.87 12.18 ;
  LAYER M2 ;
        RECT 4.57 12.04 4.89 12.32 ;
  LAYER M3 ;
        RECT 4.59 7.375 4.87 7.745 ;
  LAYER M2 ;
        RECT 4.73 7.42 6.02 7.7 ;
  LAYER M1 ;
        RECT 5.895 7.14 6.145 7.56 ;
  LAYER M2 ;
        RECT 6.02 7 7.31 7.28 ;
  LAYER M2 ;
        RECT 7.15 7 7.47 7.28 ;
  LAYER M3 ;
        RECT 7.17 7.14 7.45 7.98 ;
  LAYER M2 ;
        RECT 7.15 7.84 7.47 8.12 ;
  LAYER M2 ;
        RECT 4.57 2.8 4.89 3.08 ;
  LAYER M3 ;
        RECT 4.59 2.78 4.87 3.1 ;
  LAYER M2 ;
        RECT 4.57 12.04 4.89 12.32 ;
  LAYER M3 ;
        RECT 4.59 12.02 4.87 12.34 ;
  LAYER M2 ;
        RECT 4.57 2.8 4.89 3.08 ;
  LAYER M3 ;
        RECT 4.59 2.78 4.87 3.1 ;
  LAYER M2 ;
        RECT 4.57 12.04 4.89 12.32 ;
  LAYER M3 ;
        RECT 4.59 12.02 4.87 12.34 ;
  LAYER M1 ;
        RECT 5.895 7.055 6.145 7.225 ;
  LAYER M2 ;
        RECT 5.85 7 6.19 7.28 ;
  LAYER M1 ;
        RECT 5.895 7.475 6.145 7.645 ;
  LAYER M2 ;
        RECT 5.85 7.42 6.19 7.7 ;
  LAYER M2 ;
        RECT 4.57 2.8 4.89 3.08 ;
  LAYER M3 ;
        RECT 4.59 2.78 4.87 3.1 ;
  LAYER M2 ;
        RECT 4.57 7.42 4.89 7.7 ;
  LAYER M3 ;
        RECT 4.59 7.4 4.87 7.72 ;
  LAYER M2 ;
        RECT 4.57 12.04 4.89 12.32 ;
  LAYER M3 ;
        RECT 4.59 12.02 4.87 12.34 ;
  LAYER M1 ;
        RECT 5.895 7.055 6.145 7.225 ;
  LAYER M2 ;
        RECT 5.85 7 6.19 7.28 ;
  LAYER M1 ;
        RECT 5.895 7.475 6.145 7.645 ;
  LAYER M2 ;
        RECT 5.85 7.42 6.19 7.7 ;
  LAYER M2 ;
        RECT 4.57 2.8 4.89 3.08 ;
  LAYER M3 ;
        RECT 4.59 2.78 4.87 3.1 ;
  LAYER M2 ;
        RECT 4.57 7.42 4.89 7.7 ;
  LAYER M3 ;
        RECT 4.59 7.4 4.87 7.72 ;
  LAYER M2 ;
        RECT 4.57 12.04 4.89 12.32 ;
  LAYER M3 ;
        RECT 4.59 12.02 4.87 12.34 ;
  LAYER M1 ;
        RECT 5.895 7.055 6.145 7.225 ;
  LAYER M2 ;
        RECT 5.85 7 6.19 7.28 ;
  LAYER M1 ;
        RECT 5.895 7.475 6.145 7.645 ;
  LAYER M2 ;
        RECT 5.85 7.42 6.19 7.7 ;
  LAYER M2 ;
        RECT 4.57 2.8 4.89 3.08 ;
  LAYER M3 ;
        RECT 4.59 2.78 4.87 3.1 ;
  LAYER M2 ;
        RECT 4.57 7.42 4.89 7.7 ;
  LAYER M3 ;
        RECT 4.59 7.4 4.87 7.72 ;
  LAYER M2 ;
        RECT 4.57 12.04 4.89 12.32 ;
  LAYER M3 ;
        RECT 4.59 12.02 4.87 12.34 ;
  LAYER M2 ;
        RECT 7.15 7 7.47 7.28 ;
  LAYER M3 ;
        RECT 7.17 6.98 7.45 7.3 ;
  LAYER M2 ;
        RECT 7.15 7.84 7.47 8.12 ;
  LAYER M3 ;
        RECT 7.17 7.82 7.45 8.14 ;
  LAYER M1 ;
        RECT 5.895 7.055 6.145 7.225 ;
  LAYER M2 ;
        RECT 5.85 7 6.19 7.28 ;
  LAYER M1 ;
        RECT 5.895 7.475 6.145 7.645 ;
  LAYER M2 ;
        RECT 5.85 7.42 6.19 7.7 ;
  LAYER M2 ;
        RECT 4.57 2.8 4.89 3.08 ;
  LAYER M3 ;
        RECT 4.59 2.78 4.87 3.1 ;
  LAYER M2 ;
        RECT 4.57 7.42 4.89 7.7 ;
  LAYER M3 ;
        RECT 4.59 7.4 4.87 7.72 ;
  LAYER M2 ;
        RECT 4.57 12.04 4.89 12.32 ;
  LAYER M3 ;
        RECT 4.59 12.02 4.87 12.34 ;
  LAYER M2 ;
        RECT 7.15 7 7.47 7.28 ;
  LAYER M3 ;
        RECT 7.17 6.98 7.45 7.3 ;
  LAYER M2 ;
        RECT 7.15 7.84 7.47 8.12 ;
  LAYER M3 ;
        RECT 7.17 7.82 7.45 8.14 ;
  LAYER M1 ;
        RECT 10.625 7.895 10.875 11.425 ;
  LAYER M1 ;
        RECT 10.625 11.675 10.875 12.685 ;
  LAYER M1 ;
        RECT 10.625 13.775 10.875 14.785 ;
  LAYER M1 ;
        RECT 11.055 7.895 11.305 11.425 ;
  LAYER M1 ;
        RECT 10.195 7.895 10.445 11.425 ;
  LAYER M1 ;
        RECT 9.765 7.895 10.015 11.425 ;
  LAYER M1 ;
        RECT 9.765 11.675 10.015 12.685 ;
  LAYER M1 ;
        RECT 9.765 13.775 10.015 14.785 ;
  LAYER M1 ;
        RECT 9.335 7.895 9.585 11.425 ;
  LAYER M1 ;
        RECT 8.905 7.895 9.155 11.425 ;
  LAYER M1 ;
        RECT 8.905 11.675 9.155 12.685 ;
  LAYER M1 ;
        RECT 8.905 13.775 9.155 14.785 ;
  LAYER M1 ;
        RECT 8.475 7.895 8.725 11.425 ;
  LAYER M1 ;
        RECT 8.045 7.895 8.295 11.425 ;
  LAYER M1 ;
        RECT 8.045 11.675 8.295 12.685 ;
  LAYER M1 ;
        RECT 8.045 13.775 8.295 14.785 ;
  LAYER M1 ;
        RECT 7.615 7.895 7.865 11.425 ;
  LAYER M1 ;
        RECT 7.185 7.895 7.435 11.425 ;
  LAYER M1 ;
        RECT 7.185 11.675 7.435 12.685 ;
  LAYER M1 ;
        RECT 7.185 13.775 7.435 14.785 ;
  LAYER M1 ;
        RECT 6.755 7.895 7.005 11.425 ;
  LAYER M2 ;
        RECT 6.71 8.26 11.35 8.54 ;
  LAYER M2 ;
        RECT 7.14 14.14 10.92 14.42 ;
  LAYER M2 ;
        RECT 7.14 7.84 10.92 8.12 ;
  LAYER M2 ;
        RECT 7.14 12.04 10.92 12.32 ;
  LAYER M3 ;
        RECT 8.46 8.24 8.74 14.44 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 11.425 ;
  LAYER M1 ;
        RECT 1.165 11.675 1.415 12.685 ;
  LAYER M1 ;
        RECT 1.165 13.775 1.415 14.785 ;
  LAYER M1 ;
        RECT 0.735 7.895 0.985 11.425 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 11.425 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 11.425 ;
  LAYER M1 ;
        RECT 2.025 11.675 2.275 12.685 ;
  LAYER M1 ;
        RECT 2.025 13.775 2.275 14.785 ;
  LAYER M1 ;
        RECT 2.455 7.895 2.705 11.425 ;
  LAYER M1 ;
        RECT 2.885 7.895 3.135 11.425 ;
  LAYER M1 ;
        RECT 2.885 11.675 3.135 12.685 ;
  LAYER M1 ;
        RECT 2.885 13.775 3.135 14.785 ;
  LAYER M1 ;
        RECT 3.315 7.895 3.565 11.425 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 11.425 ;
  LAYER M1 ;
        RECT 3.745 11.675 3.995 12.685 ;
  LAYER M1 ;
        RECT 3.745 13.775 3.995 14.785 ;
  LAYER M1 ;
        RECT 4.175 7.895 4.425 11.425 ;
  LAYER M1 ;
        RECT 4.605 7.895 4.855 11.425 ;
  LAYER M1 ;
        RECT 4.605 11.675 4.855 12.685 ;
  LAYER M1 ;
        RECT 4.605 13.775 4.855 14.785 ;
  LAYER M1 ;
        RECT 5.035 7.895 5.285 11.425 ;
  LAYER M2 ;
        RECT 0.69 8.26 5.33 8.54 ;
  LAYER M2 ;
        RECT 1.12 14.14 4.9 14.42 ;
  LAYER M2 ;
        RECT 1.12 7.84 4.9 8.12 ;
  LAYER M2 ;
        RECT 1.12 12.04 4.9 12.32 ;
  LAYER M3 ;
        RECT 3.3 8.24 3.58 14.44 ;
  LAYER M1 ;
        RECT 10.625 3.695 10.875 7.225 ;
  LAYER M1 ;
        RECT 10.625 2.435 10.875 3.445 ;
  LAYER M1 ;
        RECT 10.625 0.335 10.875 1.345 ;
  LAYER M1 ;
        RECT 11.055 3.695 11.305 7.225 ;
  LAYER M1 ;
        RECT 10.195 3.695 10.445 7.225 ;
  LAYER M1 ;
        RECT 9.765 3.695 10.015 7.225 ;
  LAYER M1 ;
        RECT 9.765 2.435 10.015 3.445 ;
  LAYER M1 ;
        RECT 9.765 0.335 10.015 1.345 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M1 ;
        RECT 8.905 3.695 9.155 7.225 ;
  LAYER M1 ;
        RECT 8.905 2.435 9.155 3.445 ;
  LAYER M1 ;
        RECT 8.905 0.335 9.155 1.345 ;
  LAYER M1 ;
        RECT 8.475 3.695 8.725 7.225 ;
  LAYER M1 ;
        RECT 8.045 3.695 8.295 7.225 ;
  LAYER M1 ;
        RECT 8.045 2.435 8.295 3.445 ;
  LAYER M1 ;
        RECT 8.045 0.335 8.295 1.345 ;
  LAYER M1 ;
        RECT 7.615 3.695 7.865 7.225 ;
  LAYER M1 ;
        RECT 7.185 3.695 7.435 7.225 ;
  LAYER M1 ;
        RECT 7.185 2.435 7.435 3.445 ;
  LAYER M1 ;
        RECT 7.185 0.335 7.435 1.345 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M2 ;
        RECT 6.71 6.58 11.35 6.86 ;
  LAYER M2 ;
        RECT 7.14 0.7 10.92 0.98 ;
  LAYER M2 ;
        RECT 7.14 7 10.92 7.28 ;
  LAYER M2 ;
        RECT 7.14 2.8 10.92 3.08 ;
  LAYER M3 ;
        RECT 8.46 0.68 8.74 6.88 ;
  LAYER M1 ;
        RECT 1.165 3.695 1.415 7.225 ;
  LAYER M1 ;
        RECT 1.165 2.435 1.415 3.445 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 1.345 ;
  LAYER M1 ;
        RECT 0.735 3.695 0.985 7.225 ;
  LAYER M1 ;
        RECT 1.595 3.695 1.845 7.225 ;
  LAYER M1 ;
        RECT 2.025 3.695 2.275 7.225 ;
  LAYER M1 ;
        RECT 2.025 2.435 2.275 3.445 ;
  LAYER M1 ;
        RECT 2.025 0.335 2.275 1.345 ;
  LAYER M1 ;
        RECT 2.455 3.695 2.705 7.225 ;
  LAYER M1 ;
        RECT 2.885 3.695 3.135 7.225 ;
  LAYER M1 ;
        RECT 2.885 2.435 3.135 3.445 ;
  LAYER M1 ;
        RECT 2.885 0.335 3.135 1.345 ;
  LAYER M1 ;
        RECT 3.315 3.695 3.565 7.225 ;
  LAYER M1 ;
        RECT 3.745 3.695 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.745 2.435 3.995 3.445 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 1.345 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M1 ;
        RECT 4.605 3.695 4.855 7.225 ;
  LAYER M1 ;
        RECT 4.605 2.435 4.855 3.445 ;
  LAYER M1 ;
        RECT 4.605 0.335 4.855 1.345 ;
  LAYER M1 ;
        RECT 5.035 3.695 5.285 7.225 ;
  LAYER M2 ;
        RECT 0.69 6.58 5.33 6.86 ;
  LAYER M2 ;
        RECT 1.12 0.7 4.9 0.98 ;
  LAYER M2 ;
        RECT 1.12 7 4.9 7.28 ;
  LAYER M2 ;
        RECT 1.12 2.8 4.9 3.08 ;
  LAYER M3 ;
        RECT 3.3 0.68 3.58 6.88 ;
  LAYER M1 ;
        RECT 7.615 23.015 7.865 26.545 ;
  LAYER M1 ;
        RECT 7.615 26.795 7.865 27.805 ;
  LAYER M1 ;
        RECT 7.615 28.895 7.865 29.905 ;
  LAYER M1 ;
        RECT 8.045 23.015 8.295 26.545 ;
  LAYER M1 ;
        RECT 7.185 23.015 7.435 26.545 ;
  LAYER M1 ;
        RECT 6.755 23.015 7.005 26.545 ;
  LAYER M1 ;
        RECT 6.755 26.795 7.005 27.805 ;
  LAYER M1 ;
        RECT 6.755 28.895 7.005 29.905 ;
  LAYER M1 ;
        RECT 6.325 23.015 6.575 26.545 ;
  LAYER M1 ;
        RECT 5.895 23.015 6.145 26.545 ;
  LAYER M1 ;
        RECT 5.895 26.795 6.145 27.805 ;
  LAYER M1 ;
        RECT 5.895 28.895 6.145 29.905 ;
  LAYER M1 ;
        RECT 5.465 23.015 5.715 26.545 ;
  LAYER M1 ;
        RECT 5.035 23.015 5.285 26.545 ;
  LAYER M1 ;
        RECT 5.035 26.795 5.285 27.805 ;
  LAYER M1 ;
        RECT 5.035 28.895 5.285 29.905 ;
  LAYER M1 ;
        RECT 4.605 23.015 4.855 26.545 ;
  LAYER M1 ;
        RECT 4.175 23.015 4.425 26.545 ;
  LAYER M1 ;
        RECT 4.175 26.795 4.425 27.805 ;
  LAYER M1 ;
        RECT 4.175 28.895 4.425 29.905 ;
  LAYER M1 ;
        RECT 3.745 23.015 3.995 26.545 ;
  LAYER M2 ;
        RECT 3.7 23.38 8.34 23.66 ;
  LAYER M2 ;
        RECT 4.13 29.26 7.91 29.54 ;
  LAYER M2 ;
        RECT 4.13 22.96 7.91 23.24 ;
  LAYER M2 ;
        RECT 4.13 27.16 7.91 27.44 ;
  LAYER M3 ;
        RECT 5.45 23.36 5.73 29.56 ;
  LAYER M1 ;
        RECT 7.615 18.815 7.865 22.345 ;
  LAYER M1 ;
        RECT 7.615 17.555 7.865 18.565 ;
  LAYER M1 ;
        RECT 7.615 15.455 7.865 16.465 ;
  LAYER M1 ;
        RECT 8.045 18.815 8.295 22.345 ;
  LAYER M1 ;
        RECT 7.185 18.815 7.435 22.345 ;
  LAYER M1 ;
        RECT 6.755 18.815 7.005 22.345 ;
  LAYER M1 ;
        RECT 6.755 17.555 7.005 18.565 ;
  LAYER M1 ;
        RECT 6.755 15.455 7.005 16.465 ;
  LAYER M1 ;
        RECT 6.325 18.815 6.575 22.345 ;
  LAYER M1 ;
        RECT 5.895 18.815 6.145 22.345 ;
  LAYER M1 ;
        RECT 5.895 17.555 6.145 18.565 ;
  LAYER M1 ;
        RECT 5.895 15.455 6.145 16.465 ;
  LAYER M1 ;
        RECT 5.465 18.815 5.715 22.345 ;
  LAYER M1 ;
        RECT 5.035 18.815 5.285 22.345 ;
  LAYER M1 ;
        RECT 5.035 17.555 5.285 18.565 ;
  LAYER M1 ;
        RECT 5.035 15.455 5.285 16.465 ;
  LAYER M1 ;
        RECT 4.605 18.815 4.855 22.345 ;
  LAYER M1 ;
        RECT 4.175 18.815 4.425 22.345 ;
  LAYER M1 ;
        RECT 4.175 17.555 4.425 18.565 ;
  LAYER M1 ;
        RECT 4.175 15.455 4.425 16.465 ;
  LAYER M1 ;
        RECT 3.745 18.815 3.995 22.345 ;
  LAYER M2 ;
        RECT 3.7 21.7 8.34 21.98 ;
  LAYER M2 ;
        RECT 4.13 15.82 7.91 16.1 ;
  LAYER M2 ;
        RECT 4.13 22.12 7.91 22.4 ;
  LAYER M2 ;
        RECT 4.13 17.92 7.91 18.2 ;
  LAYER M3 ;
        RECT 5.45 15.8 5.73 22 ;
  END 
END RINGOSC
