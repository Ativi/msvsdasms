module ONEBITADC_0(
     input Vin,
     input vref,
     output out
);

endmodule
