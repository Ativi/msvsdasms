VERSION 5.7 ;

  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO STAGE2_INV_62673116_0_0_1679063325
  CLASS BLOCK ;
  FOREIGN STAGE2_INV_62673116_0_0_1679063325 ;
  ORIGIN 0.000 -0.150 ;
  SIZE 12.040 BY 14.970 ;
  OBS
      LAYER nwell ;
        RECT 0.000 7.560 12.040 15.120 ;
      LAYER pwell ;
        RECT 0.605 4.070 5.415 5.380 ;
        RECT 6.625 4.070 11.435 5.380 ;
        RECT 1.075 0.150 4.945 1.530 ;
        RECT 7.095 0.150 10.965 1.530 ;
      LAYER li1 ;
        RECT 1.165 13.775 1.415 14.785 ;
        RECT 2.025 13.775 2.275 14.785 ;
        RECT 2.885 13.775 3.135 14.785 ;
        RECT 3.745 13.775 3.995 14.785 ;
        RECT 4.605 13.775 4.855 14.785 ;
        RECT 7.185 13.775 7.435 14.785 ;
        RECT 8.045 13.775 8.295 14.785 ;
        RECT 8.905 13.775 9.155 14.785 ;
        RECT 9.765 13.775 10.015 14.785 ;
        RECT 10.625 13.775 10.875 14.785 ;
        RECT 1.165 11.675 1.415 12.685 ;
        RECT 2.025 11.675 2.275 12.685 ;
        RECT 2.885 11.675 3.135 12.685 ;
        RECT 3.745 11.675 3.995 12.685 ;
        RECT 4.605 11.675 4.855 12.685 ;
        RECT 7.185 11.675 7.435 12.685 ;
        RECT 8.045 11.675 8.295 12.685 ;
        RECT 8.905 11.675 9.155 12.685 ;
        RECT 9.765 11.675 10.015 12.685 ;
        RECT 10.625 11.675 10.875 12.685 ;
        RECT 0.735 7.895 0.985 11.425 ;
        RECT 1.165 7.895 1.415 11.425 ;
        RECT 1.595 7.895 1.845 11.425 ;
        RECT 2.025 7.895 2.275 11.425 ;
        RECT 2.455 7.895 2.705 11.425 ;
        RECT 2.885 7.895 3.135 11.425 ;
        RECT 3.315 7.895 3.565 11.425 ;
        RECT 3.745 7.895 3.995 11.425 ;
        RECT 4.175 7.895 4.425 11.425 ;
        RECT 4.605 7.895 4.855 11.425 ;
        RECT 5.035 7.895 5.285 11.425 ;
        RECT 5.895 7.475 6.145 8.065 ;
        RECT 6.755 7.895 7.005 11.425 ;
        RECT 7.185 7.895 7.435 11.425 ;
        RECT 7.615 7.895 7.865 11.425 ;
        RECT 8.045 7.895 8.295 11.425 ;
        RECT 8.475 7.895 8.725 11.425 ;
        RECT 8.905 7.895 9.155 11.425 ;
        RECT 9.335 7.895 9.585 11.425 ;
        RECT 9.765 7.895 10.015 11.425 ;
        RECT 10.195 7.895 10.445 11.425 ;
        RECT 10.625 7.895 10.875 11.425 ;
        RECT 11.055 7.895 11.305 11.425 ;
        RECT 0.735 3.695 0.985 7.225 ;
        RECT 1.165 3.695 1.415 7.225 ;
        RECT 1.595 3.695 1.845 7.225 ;
        RECT 2.025 3.695 2.275 7.225 ;
        RECT 2.455 3.695 2.705 7.225 ;
        RECT 2.885 3.695 3.135 7.225 ;
        RECT 3.315 3.695 3.565 7.225 ;
        RECT 3.745 3.695 3.995 7.225 ;
        RECT 4.175 3.695 4.425 7.225 ;
        RECT 4.605 3.695 4.855 7.225 ;
        RECT 5.035 3.695 5.285 7.225 ;
        RECT 6.755 3.695 7.005 7.225 ;
        RECT 7.185 3.695 7.435 7.225 ;
        RECT 7.615 3.695 7.865 7.225 ;
        RECT 8.045 3.695 8.295 7.225 ;
        RECT 8.475 3.695 8.725 7.225 ;
        RECT 8.905 3.695 9.155 7.225 ;
        RECT 9.335 3.695 9.585 7.225 ;
        RECT 9.765 3.695 10.015 7.225 ;
        RECT 10.195 3.695 10.445 7.225 ;
        RECT 10.625 3.695 10.875 7.225 ;
        RECT 11.055 3.695 11.305 7.225 ;
        RECT 1.165 2.435 1.415 3.445 ;
        RECT 2.025 2.435 2.275 3.445 ;
        RECT 2.885 2.435 3.135 3.445 ;
        RECT 3.745 2.435 3.995 3.445 ;
        RECT 4.605 2.435 4.855 3.445 ;
        RECT 7.185 2.435 7.435 3.445 ;
        RECT 8.045 2.435 8.295 3.445 ;
        RECT 8.905 2.435 9.155 3.445 ;
        RECT 9.765 2.435 10.015 3.445 ;
        RECT 10.625 2.435 10.875 3.445 ;
        RECT 1.165 0.335 1.415 1.345 ;
        RECT 2.025 0.335 2.275 1.345 ;
        RECT 2.885 0.335 3.135 1.345 ;
        RECT 3.745 0.335 3.995 1.345 ;
        RECT 4.605 0.335 4.855 1.345 ;
        RECT 7.185 0.335 7.435 1.345 ;
        RECT 8.045 0.335 8.295 1.345 ;
        RECT 8.905 0.335 9.155 1.345 ;
        RECT 9.765 0.335 10.015 1.345 ;
        RECT 10.625 0.335 10.875 1.345 ;
      LAYER mcon ;
        RECT 1.205 14.195 1.375 14.365 ;
        RECT 2.065 14.195 2.235 14.365 ;
        RECT 2.925 14.195 3.095 14.365 ;
        RECT 3.785 14.195 3.955 14.365 ;
        RECT 4.645 14.195 4.815 14.365 ;
        RECT 7.225 14.195 7.395 14.365 ;
        RECT 8.085 14.195 8.255 14.365 ;
        RECT 8.945 14.195 9.115 14.365 ;
        RECT 9.805 14.195 9.975 14.365 ;
        RECT 10.665 14.195 10.835 14.365 ;
        RECT 1.205 12.095 1.375 12.265 ;
        RECT 2.065 12.095 2.235 12.265 ;
        RECT 2.925 12.095 3.095 12.265 ;
        RECT 3.785 12.095 3.955 12.265 ;
        RECT 4.645 12.095 4.815 12.265 ;
        RECT 7.225 12.095 7.395 12.265 ;
        RECT 8.085 12.095 8.255 12.265 ;
        RECT 8.945 12.095 9.115 12.265 ;
        RECT 9.805 12.095 9.975 12.265 ;
        RECT 10.665 12.095 10.835 12.265 ;
        RECT 0.775 8.315 0.945 8.485 ;
        RECT 1.205 7.895 1.375 8.065 ;
        RECT 1.635 8.315 1.805 8.485 ;
        RECT 2.065 7.895 2.235 8.065 ;
        RECT 2.495 8.315 2.665 8.485 ;
        RECT 2.925 7.895 3.095 8.065 ;
        RECT 3.355 8.315 3.525 8.485 ;
        RECT 3.785 7.895 3.955 8.065 ;
        RECT 4.215 8.315 4.385 8.485 ;
        RECT 4.645 7.895 4.815 8.065 ;
        RECT 5.075 8.315 5.245 8.485 ;
        RECT 6.795 8.315 6.965 8.485 ;
        RECT 5.935 7.895 6.105 8.065 ;
        RECT 7.225 7.895 7.395 8.065 ;
        RECT 7.655 8.315 7.825 8.485 ;
        RECT 8.085 7.895 8.255 8.065 ;
        RECT 8.515 8.315 8.685 8.485 ;
        RECT 8.945 7.895 9.115 8.065 ;
        RECT 9.375 8.315 9.545 8.485 ;
        RECT 9.805 7.895 9.975 8.065 ;
        RECT 10.235 8.315 10.405 8.485 ;
        RECT 10.665 7.895 10.835 8.065 ;
        RECT 11.095 8.315 11.265 8.485 ;
        RECT 5.935 7.475 6.105 7.645 ;
        RECT 0.775 6.635 0.945 6.805 ;
        RECT 1.205 7.055 1.375 7.225 ;
        RECT 1.635 6.635 1.805 6.805 ;
        RECT 2.065 7.055 2.235 7.225 ;
        RECT 2.495 6.635 2.665 6.805 ;
        RECT 2.925 7.055 3.095 7.225 ;
        RECT 3.355 6.635 3.525 6.805 ;
        RECT 3.785 7.055 3.955 7.225 ;
        RECT 4.215 6.635 4.385 6.805 ;
        RECT 4.645 7.055 4.815 7.225 ;
        RECT 5.075 6.635 5.245 6.805 ;
        RECT 6.795 6.635 6.965 6.805 ;
        RECT 7.225 7.055 7.395 7.225 ;
        RECT 7.655 6.635 7.825 6.805 ;
        RECT 8.085 7.055 8.255 7.225 ;
        RECT 8.515 6.635 8.685 6.805 ;
        RECT 8.945 7.055 9.115 7.225 ;
        RECT 9.375 6.635 9.545 6.805 ;
        RECT 9.805 7.055 9.975 7.225 ;
        RECT 10.235 6.635 10.405 6.805 ;
        RECT 10.665 7.055 10.835 7.225 ;
        RECT 11.095 6.635 11.265 6.805 ;
        RECT 1.205 2.855 1.375 3.025 ;
        RECT 2.065 2.855 2.235 3.025 ;
        RECT 2.925 2.855 3.095 3.025 ;
        RECT 3.785 2.855 3.955 3.025 ;
        RECT 4.645 2.855 4.815 3.025 ;
        RECT 7.225 2.855 7.395 3.025 ;
        RECT 8.085 2.855 8.255 3.025 ;
        RECT 8.945 2.855 9.115 3.025 ;
        RECT 9.805 2.855 9.975 3.025 ;
        RECT 10.665 2.855 10.835 3.025 ;
        RECT 1.205 0.755 1.375 0.925 ;
        RECT 2.065 0.755 2.235 0.925 ;
        RECT 2.925 0.755 3.095 0.925 ;
        RECT 3.785 0.755 3.955 0.925 ;
        RECT 4.645 0.755 4.815 0.925 ;
        RECT 7.225 0.755 7.395 0.925 ;
        RECT 8.085 0.755 8.255 0.925 ;
        RECT 8.945 0.755 9.115 0.925 ;
        RECT 9.805 0.755 9.975 0.925 ;
        RECT 10.665 0.755 10.835 0.925 ;
      LAYER met1 ;
        RECT 1.120 14.140 4.900 14.420 ;
        RECT 7.140 14.140 10.920 14.420 ;
        RECT 1.120 12.040 4.900 12.320 ;
        RECT 7.140 12.040 10.920 12.320 ;
        RECT 3.280 11.200 8.760 11.480 ;
        RECT 0.690 8.260 5.330 8.540 ;
        RECT 6.710 8.260 11.350 8.540 ;
        RECT 1.120 7.840 4.900 8.120 ;
        RECT 5.850 7.840 10.920 8.120 ;
        RECT 4.570 7.420 6.190 7.700 ;
        RECT 1.120 7.000 4.900 7.280 ;
        RECT 7.140 7.000 10.920 7.280 ;
        RECT 0.690 6.580 5.330 6.860 ;
        RECT 6.710 6.580 11.350 6.860 ;
        RECT 3.280 3.640 8.760 3.920 ;
        RECT 1.120 2.800 4.900 3.080 ;
        RECT 7.140 2.800 10.920 3.080 ;
        RECT 1.120 0.700 4.900 0.980 ;
        RECT 7.140 0.700 10.920 0.980 ;
      LAYER via ;
        RECT 3.310 14.150 3.570 14.410 ;
        RECT 8.470 14.150 8.730 14.410 ;
        RECT 4.600 12.050 4.860 12.310 ;
        RECT 8.900 12.050 9.160 12.310 ;
        RECT 3.310 11.210 3.570 11.470 ;
        RECT 8.470 11.210 8.730 11.470 ;
        RECT 3.310 8.270 3.570 8.530 ;
        RECT 8.470 8.270 8.730 8.530 ;
        RECT 2.880 7.850 3.140 8.110 ;
        RECT 7.180 7.850 7.440 8.110 ;
        RECT 4.600 7.430 4.860 7.690 ;
        RECT 2.880 7.010 3.140 7.270 ;
        RECT 7.180 7.010 7.440 7.270 ;
        RECT 3.310 6.590 3.570 6.850 ;
        RECT 8.470 6.590 8.730 6.850 ;
        RECT 3.310 3.650 3.570 3.910 ;
        RECT 8.470 3.650 8.730 3.910 ;
        RECT 4.600 2.810 4.860 3.070 ;
        RECT 8.900 2.810 9.160 3.070 ;
        RECT 3.310 0.710 3.570 0.970 ;
        RECT 8.470 0.710 8.730 0.970 ;
      LAYER met2 ;
        RECT 3.300 8.240 3.580 14.440 ;
        RECT 2.870 6.980 3.150 8.140 ;
        RECT 3.300 0.680 3.580 6.880 ;
        RECT 4.590 2.780 4.870 12.340 ;
        RECT 8.460 8.240 8.740 14.440 ;
        RECT 7.170 6.980 7.450 8.140 ;
        RECT 8.460 0.680 8.740 6.880 ;
        RECT 8.890 2.780 9.170 12.340 ;
  END
END STAGE2_INV_62673116_0_0_1679063325
MACRO INV_57920576_0_0_1679063324
  CLASS BLOCK ;
  FOREIGN INV_57920576_0_0_1679063324 ;
  ORIGIN 0.000 -0.150 ;
  SIZE 6.020 BY 14.970 ;
  OBS
      LAYER nwell ;
        RECT 0.000 7.560 6.020 15.120 ;
      LAYER pwell ;
        RECT 0.605 4.070 5.415 5.380 ;
        RECT 1.075 0.150 4.945 1.530 ;
      LAYER li1 ;
        RECT 1.165 13.775 1.415 14.785 ;
        RECT 2.025 13.775 2.275 14.785 ;
        RECT 2.885 13.775 3.135 14.785 ;
        RECT 3.745 13.775 3.995 14.785 ;
        RECT 4.605 13.775 4.855 14.785 ;
        RECT 1.165 11.675 1.415 12.685 ;
        RECT 2.025 11.675 2.275 12.685 ;
        RECT 2.885 11.675 3.135 12.685 ;
        RECT 3.745 11.675 3.995 12.685 ;
        RECT 4.605 11.675 4.855 12.685 ;
        RECT 0.735 7.895 0.985 11.425 ;
        RECT 1.165 7.895 1.415 11.425 ;
        RECT 1.595 7.895 1.845 11.425 ;
        RECT 2.025 7.895 2.275 11.425 ;
        RECT 2.455 7.895 2.705 11.425 ;
        RECT 2.885 7.895 3.135 11.425 ;
        RECT 3.315 7.895 3.565 11.425 ;
        RECT 3.745 7.895 3.995 11.425 ;
        RECT 4.175 7.895 4.425 11.425 ;
        RECT 4.605 7.895 4.855 11.425 ;
        RECT 5.035 7.895 5.285 11.425 ;
        RECT 0.735 3.695 0.985 7.225 ;
        RECT 1.165 3.695 1.415 7.225 ;
        RECT 1.595 3.695 1.845 7.225 ;
        RECT 2.025 3.695 2.275 7.225 ;
        RECT 2.455 3.695 2.705 7.225 ;
        RECT 2.885 3.695 3.135 7.225 ;
        RECT 3.315 3.695 3.565 7.225 ;
        RECT 3.745 3.695 3.995 7.225 ;
        RECT 4.175 3.695 4.425 7.225 ;
        RECT 4.605 3.695 4.855 7.225 ;
        RECT 5.035 3.695 5.285 7.225 ;
        RECT 1.165 2.435 1.415 3.445 ;
        RECT 2.025 2.435 2.275 3.445 ;
        RECT 2.885 2.435 3.135 3.445 ;
        RECT 3.745 2.435 3.995 3.445 ;
        RECT 4.605 2.435 4.855 3.445 ;
        RECT 1.165 0.335 1.415 1.345 ;
        RECT 2.025 0.335 2.275 1.345 ;
        RECT 2.885 0.335 3.135 1.345 ;
        RECT 3.745 0.335 3.995 1.345 ;
        RECT 4.605 0.335 4.855 1.345 ;
      LAYER mcon ;
        RECT 1.205 14.195 1.375 14.365 ;
        RECT 2.065 14.195 2.235 14.365 ;
        RECT 2.925 14.195 3.095 14.365 ;
        RECT 3.785 14.195 3.955 14.365 ;
        RECT 4.645 14.195 4.815 14.365 ;
        RECT 1.205 12.095 1.375 12.265 ;
        RECT 2.065 12.095 2.235 12.265 ;
        RECT 2.925 12.095 3.095 12.265 ;
        RECT 3.785 12.095 3.955 12.265 ;
        RECT 4.645 12.095 4.815 12.265 ;
        RECT 0.775 8.315 0.945 8.485 ;
        RECT 1.205 7.895 1.375 8.065 ;
        RECT 1.635 8.315 1.805 8.485 ;
        RECT 2.065 7.895 2.235 8.065 ;
        RECT 2.495 8.315 2.665 8.485 ;
        RECT 2.925 7.895 3.095 8.065 ;
        RECT 3.355 8.315 3.525 8.485 ;
        RECT 3.785 7.895 3.955 8.065 ;
        RECT 4.215 8.315 4.385 8.485 ;
        RECT 4.645 7.895 4.815 8.065 ;
        RECT 5.075 8.315 5.245 8.485 ;
        RECT 0.775 6.635 0.945 6.805 ;
        RECT 1.205 7.055 1.375 7.225 ;
        RECT 1.635 6.635 1.805 6.805 ;
        RECT 2.065 7.055 2.235 7.225 ;
        RECT 2.495 6.635 2.665 6.805 ;
        RECT 2.925 7.055 3.095 7.225 ;
        RECT 3.355 6.635 3.525 6.805 ;
        RECT 3.785 7.055 3.955 7.225 ;
        RECT 4.215 6.635 4.385 6.805 ;
        RECT 4.645 7.055 4.815 7.225 ;
        RECT 5.075 6.635 5.245 6.805 ;
        RECT 1.205 2.855 1.375 3.025 ;
        RECT 2.065 2.855 2.235 3.025 ;
        RECT 2.925 2.855 3.095 3.025 ;
        RECT 3.785 2.855 3.955 3.025 ;
        RECT 4.645 2.855 4.815 3.025 ;
        RECT 1.205 0.755 1.375 0.925 ;
        RECT 2.065 0.755 2.235 0.925 ;
        RECT 2.925 0.755 3.095 0.925 ;
        RECT 3.785 0.755 3.955 0.925 ;
        RECT 4.645 0.755 4.815 0.925 ;
      LAYER met1 ;
        RECT 1.120 14.140 4.900 14.420 ;
        RECT 1.120 12.040 4.900 12.320 ;
        RECT 0.690 8.260 5.330 8.540 ;
        RECT 1.120 7.840 4.900 8.120 ;
        RECT 1.120 7.000 4.900 7.280 ;
        RECT 0.690 6.580 5.330 6.860 ;
        RECT 1.120 2.800 4.900 3.080 ;
        RECT 1.120 0.700 4.900 0.980 ;
      LAYER via ;
        RECT 2.450 14.150 2.710 14.410 ;
        RECT 3.310 12.050 3.570 12.310 ;
        RECT 2.450 8.270 2.710 8.530 ;
        RECT 2.880 7.850 3.140 8.110 ;
        RECT 2.880 7.010 3.140 7.270 ;
        RECT 2.450 6.590 2.710 6.850 ;
        RECT 3.310 2.810 3.570 3.070 ;
        RECT 2.450 0.710 2.710 0.970 ;
      LAYER met2 ;
        RECT 2.440 8.240 2.720 14.440 ;
        RECT 2.870 6.980 3.150 8.140 ;
        RECT 2.440 0.680 2.720 6.880 ;
        RECT 3.300 2.780 3.580 12.340 ;
  END
END INV_57920576_0_0_1679063324
MACRO RINGOSC_0
  CLASS BLOCK ;
  FOREIGN RINGOSC_0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.040 BY 30.090 ;
  OBS
      LAYER pwell ;
        RECT 4.085 28.710 7.955 30.090 ;
        RECT 3.615 24.860 8.425 26.170 ;
      LAYER nwell ;
        RECT 3.010 15.120 9.030 22.680 ;
      LAYER pwell ;
        RECT 1.075 13.590 4.945 14.970 ;
        RECT 7.095 13.590 10.965 14.970 ;
        RECT 0.605 9.740 5.415 11.050 ;
        RECT 6.625 9.740 11.435 11.050 ;
      LAYER nwell ;
        RECT 0.000 0.000 12.040 7.560 ;
      LAYER li1 ;
        RECT 4.175 28.895 4.425 29.905 ;
        RECT 5.035 28.895 5.285 29.905 ;
        RECT 5.895 28.895 6.145 29.905 ;
        RECT 6.755 28.895 7.005 29.905 ;
        RECT 7.615 28.895 7.865 29.905 ;
        RECT 4.175 26.795 4.425 27.805 ;
        RECT 5.035 26.795 5.285 27.805 ;
        RECT 5.895 26.795 6.145 27.805 ;
        RECT 6.755 26.795 7.005 27.805 ;
        RECT 7.615 26.795 7.865 27.805 ;
        RECT 3.745 23.015 3.995 26.545 ;
        RECT 4.175 23.015 4.425 26.545 ;
        RECT 4.605 23.015 4.855 26.545 ;
        RECT 5.035 23.015 5.285 26.545 ;
        RECT 5.465 23.015 5.715 26.545 ;
        RECT 5.895 23.015 6.145 26.545 ;
        RECT 6.325 23.015 6.575 26.545 ;
        RECT 6.755 23.015 7.005 26.545 ;
        RECT 7.185 23.015 7.435 26.545 ;
        RECT 7.615 23.015 7.865 26.545 ;
        RECT 8.045 23.015 8.295 26.545 ;
        RECT 3.745 18.815 3.995 22.345 ;
        RECT 4.175 18.815 4.425 22.345 ;
        RECT 4.605 18.815 4.855 22.345 ;
        RECT 5.035 18.815 5.285 22.345 ;
        RECT 5.465 18.815 5.715 22.345 ;
        RECT 5.895 18.815 6.145 22.345 ;
        RECT 6.325 18.815 6.575 22.345 ;
        RECT 6.755 18.815 7.005 22.345 ;
        RECT 7.185 18.815 7.435 22.345 ;
        RECT 7.615 18.815 7.865 22.345 ;
        RECT 8.045 18.815 8.295 22.345 ;
        RECT 4.175 17.555 4.425 18.565 ;
        RECT 5.035 17.555 5.285 18.565 ;
        RECT 5.895 17.555 6.145 18.565 ;
        RECT 6.755 17.555 7.005 18.565 ;
        RECT 7.615 17.555 7.865 18.565 ;
        RECT 4.175 15.455 4.425 16.465 ;
        RECT 5.035 15.455 5.285 16.465 ;
        RECT 5.895 15.455 6.145 16.465 ;
        RECT 6.755 15.455 7.005 16.465 ;
        RECT 7.615 15.455 7.865 16.465 ;
        RECT 1.165 13.775 1.415 14.785 ;
        RECT 2.025 13.775 2.275 14.785 ;
        RECT 2.885 13.775 3.135 14.785 ;
        RECT 3.745 13.775 3.995 14.785 ;
        RECT 4.605 13.775 4.855 14.785 ;
        RECT 7.185 13.775 7.435 14.785 ;
        RECT 8.045 13.775 8.295 14.785 ;
        RECT 8.905 13.775 9.155 14.785 ;
        RECT 9.765 13.775 10.015 14.785 ;
        RECT 10.625 13.775 10.875 14.785 ;
        RECT 1.165 11.675 1.415 12.685 ;
        RECT 2.025 11.675 2.275 12.685 ;
        RECT 2.885 11.675 3.135 12.685 ;
        RECT 3.745 11.675 3.995 12.685 ;
        RECT 4.605 11.675 4.855 12.685 ;
        RECT 7.185 11.675 7.435 12.685 ;
        RECT 8.045 11.675 8.295 12.685 ;
        RECT 8.905 11.675 9.155 12.685 ;
        RECT 9.765 11.675 10.015 12.685 ;
        RECT 10.625 11.675 10.875 12.685 ;
        RECT 0.735 7.895 0.985 11.425 ;
        RECT 1.165 7.895 1.415 11.425 ;
        RECT 1.595 7.895 1.845 11.425 ;
        RECT 2.025 7.895 2.275 11.425 ;
        RECT 2.455 7.895 2.705 11.425 ;
        RECT 2.885 7.895 3.135 11.425 ;
        RECT 3.315 7.895 3.565 11.425 ;
        RECT 3.745 7.895 3.995 11.425 ;
        RECT 4.175 7.895 4.425 11.425 ;
        RECT 4.605 7.895 4.855 11.425 ;
        RECT 5.035 7.895 5.285 11.425 ;
        RECT 6.755 7.895 7.005 11.425 ;
        RECT 7.185 7.895 7.435 11.425 ;
        RECT 7.615 7.895 7.865 11.425 ;
        RECT 8.045 7.895 8.295 11.425 ;
        RECT 8.475 7.895 8.725 11.425 ;
        RECT 8.905 7.895 9.155 11.425 ;
        RECT 9.335 7.895 9.585 11.425 ;
        RECT 9.765 7.895 10.015 11.425 ;
        RECT 10.195 7.895 10.445 11.425 ;
        RECT 10.625 7.895 10.875 11.425 ;
        RECT 11.055 7.895 11.305 11.425 ;
        RECT 0.735 3.695 0.985 7.225 ;
        RECT 1.165 3.695 1.415 7.225 ;
        RECT 1.595 3.695 1.845 7.225 ;
        RECT 2.025 3.695 2.275 7.225 ;
        RECT 2.455 3.695 2.705 7.225 ;
        RECT 2.885 3.695 3.135 7.225 ;
        RECT 3.315 3.695 3.565 7.225 ;
        RECT 3.745 3.695 3.995 7.225 ;
        RECT 4.175 3.695 4.425 7.225 ;
        RECT 4.605 3.695 4.855 7.225 ;
        RECT 5.035 3.695 5.285 7.225 ;
        RECT 5.895 7.055 6.145 7.645 ;
        RECT 6.755 3.695 7.005 7.225 ;
        RECT 7.185 3.695 7.435 7.225 ;
        RECT 7.615 3.695 7.865 7.225 ;
        RECT 8.045 3.695 8.295 7.225 ;
        RECT 8.475 3.695 8.725 7.225 ;
        RECT 8.905 3.695 9.155 7.225 ;
        RECT 9.335 3.695 9.585 7.225 ;
        RECT 9.765 3.695 10.015 7.225 ;
        RECT 10.195 3.695 10.445 7.225 ;
        RECT 10.625 3.695 10.875 7.225 ;
        RECT 11.055 3.695 11.305 7.225 ;
        RECT 1.165 2.435 1.415 3.445 ;
        RECT 2.025 2.435 2.275 3.445 ;
        RECT 2.885 2.435 3.135 3.445 ;
        RECT 3.745 2.435 3.995 3.445 ;
        RECT 4.605 2.435 4.855 3.445 ;
        RECT 7.185 2.435 7.435 3.445 ;
        RECT 8.045 2.435 8.295 3.445 ;
        RECT 8.905 2.435 9.155 3.445 ;
        RECT 9.765 2.435 10.015 3.445 ;
        RECT 10.625 2.435 10.875 3.445 ;
        RECT 1.165 0.335 1.415 1.345 ;
        RECT 2.025 0.335 2.275 1.345 ;
        RECT 2.885 0.335 3.135 1.345 ;
        RECT 3.745 0.335 3.995 1.345 ;
        RECT 4.605 0.335 4.855 1.345 ;
        RECT 7.185 0.335 7.435 1.345 ;
        RECT 8.045 0.335 8.295 1.345 ;
        RECT 8.905 0.335 9.155 1.345 ;
        RECT 9.765 0.335 10.015 1.345 ;
        RECT 10.625 0.335 10.875 1.345 ;
      LAYER mcon ;
        RECT 4.215 29.315 4.385 29.485 ;
        RECT 5.075 29.315 5.245 29.485 ;
        RECT 5.935 29.315 6.105 29.485 ;
        RECT 6.795 29.315 6.965 29.485 ;
        RECT 7.655 29.315 7.825 29.485 ;
        RECT 4.215 27.215 4.385 27.385 ;
        RECT 5.075 27.215 5.245 27.385 ;
        RECT 5.935 27.215 6.105 27.385 ;
        RECT 6.795 27.215 6.965 27.385 ;
        RECT 7.655 27.215 7.825 27.385 ;
        RECT 3.785 23.435 3.955 23.605 ;
        RECT 4.215 23.015 4.385 23.185 ;
        RECT 4.645 23.435 4.815 23.605 ;
        RECT 5.075 23.015 5.245 23.185 ;
        RECT 5.505 23.435 5.675 23.605 ;
        RECT 5.935 23.015 6.105 23.185 ;
        RECT 6.365 23.435 6.535 23.605 ;
        RECT 6.795 23.015 6.965 23.185 ;
        RECT 7.225 23.435 7.395 23.605 ;
        RECT 7.655 23.015 7.825 23.185 ;
        RECT 8.085 23.435 8.255 23.605 ;
        RECT 3.785 21.755 3.955 21.925 ;
        RECT 4.215 22.175 4.385 22.345 ;
        RECT 4.645 21.755 4.815 21.925 ;
        RECT 5.075 22.175 5.245 22.345 ;
        RECT 5.505 21.755 5.675 21.925 ;
        RECT 5.935 22.175 6.105 22.345 ;
        RECT 6.365 21.755 6.535 21.925 ;
        RECT 6.795 22.175 6.965 22.345 ;
        RECT 7.225 21.755 7.395 21.925 ;
        RECT 7.655 22.175 7.825 22.345 ;
        RECT 8.085 21.755 8.255 21.925 ;
        RECT 4.215 17.975 4.385 18.145 ;
        RECT 5.075 17.975 5.245 18.145 ;
        RECT 5.935 17.975 6.105 18.145 ;
        RECT 6.795 17.975 6.965 18.145 ;
        RECT 7.655 17.975 7.825 18.145 ;
        RECT 4.215 15.875 4.385 16.045 ;
        RECT 5.075 15.875 5.245 16.045 ;
        RECT 5.935 15.875 6.105 16.045 ;
        RECT 6.795 15.875 6.965 16.045 ;
        RECT 7.655 15.875 7.825 16.045 ;
        RECT 1.205 14.195 1.375 14.365 ;
        RECT 2.065 14.195 2.235 14.365 ;
        RECT 2.925 14.195 3.095 14.365 ;
        RECT 3.785 14.195 3.955 14.365 ;
        RECT 4.645 14.195 4.815 14.365 ;
        RECT 7.225 14.195 7.395 14.365 ;
        RECT 8.085 14.195 8.255 14.365 ;
        RECT 8.945 14.195 9.115 14.365 ;
        RECT 9.805 14.195 9.975 14.365 ;
        RECT 10.665 14.195 10.835 14.365 ;
        RECT 1.205 12.095 1.375 12.265 ;
        RECT 2.065 12.095 2.235 12.265 ;
        RECT 2.925 12.095 3.095 12.265 ;
        RECT 3.785 12.095 3.955 12.265 ;
        RECT 4.645 12.095 4.815 12.265 ;
        RECT 7.225 12.095 7.395 12.265 ;
        RECT 8.085 12.095 8.255 12.265 ;
        RECT 8.945 12.095 9.115 12.265 ;
        RECT 9.805 12.095 9.975 12.265 ;
        RECT 10.665 12.095 10.835 12.265 ;
        RECT 0.775 8.315 0.945 8.485 ;
        RECT 1.205 7.895 1.375 8.065 ;
        RECT 1.635 8.315 1.805 8.485 ;
        RECT 2.065 7.895 2.235 8.065 ;
        RECT 2.495 8.315 2.665 8.485 ;
        RECT 2.925 7.895 3.095 8.065 ;
        RECT 3.355 8.315 3.525 8.485 ;
        RECT 3.785 7.895 3.955 8.065 ;
        RECT 4.215 8.315 4.385 8.485 ;
        RECT 4.645 7.895 4.815 8.065 ;
        RECT 5.075 8.315 5.245 8.485 ;
        RECT 6.795 8.315 6.965 8.485 ;
        RECT 7.225 7.895 7.395 8.065 ;
        RECT 7.655 8.315 7.825 8.485 ;
        RECT 8.085 7.895 8.255 8.065 ;
        RECT 8.515 8.315 8.685 8.485 ;
        RECT 8.945 7.895 9.115 8.065 ;
        RECT 9.375 8.315 9.545 8.485 ;
        RECT 9.805 7.895 9.975 8.065 ;
        RECT 10.235 8.315 10.405 8.485 ;
        RECT 10.665 7.895 10.835 8.065 ;
        RECT 11.095 8.315 11.265 8.485 ;
        RECT 5.935 7.475 6.105 7.645 ;
        RECT 0.775 6.635 0.945 6.805 ;
        RECT 1.205 7.055 1.375 7.225 ;
        RECT 1.635 6.635 1.805 6.805 ;
        RECT 2.065 7.055 2.235 7.225 ;
        RECT 2.495 6.635 2.665 6.805 ;
        RECT 2.925 7.055 3.095 7.225 ;
        RECT 3.355 6.635 3.525 6.805 ;
        RECT 3.785 7.055 3.955 7.225 ;
        RECT 4.215 6.635 4.385 6.805 ;
        RECT 4.645 7.055 4.815 7.225 ;
        RECT 5.935 7.055 6.105 7.225 ;
        RECT 5.075 6.635 5.245 6.805 ;
        RECT 6.795 6.635 6.965 6.805 ;
        RECT 7.225 7.055 7.395 7.225 ;
        RECT 7.655 6.635 7.825 6.805 ;
        RECT 8.085 7.055 8.255 7.225 ;
        RECT 8.515 6.635 8.685 6.805 ;
        RECT 8.945 7.055 9.115 7.225 ;
        RECT 9.375 6.635 9.545 6.805 ;
        RECT 9.805 7.055 9.975 7.225 ;
        RECT 10.235 6.635 10.405 6.805 ;
        RECT 10.665 7.055 10.835 7.225 ;
        RECT 11.095 6.635 11.265 6.805 ;
        RECT 1.205 2.855 1.375 3.025 ;
        RECT 2.065 2.855 2.235 3.025 ;
        RECT 2.925 2.855 3.095 3.025 ;
        RECT 3.785 2.855 3.955 3.025 ;
        RECT 4.645 2.855 4.815 3.025 ;
        RECT 7.225 2.855 7.395 3.025 ;
        RECT 8.085 2.855 8.255 3.025 ;
        RECT 8.945 2.855 9.115 3.025 ;
        RECT 9.805 2.855 9.975 3.025 ;
        RECT 10.665 2.855 10.835 3.025 ;
        RECT 1.205 0.755 1.375 0.925 ;
        RECT 2.065 0.755 2.235 0.925 ;
        RECT 2.925 0.755 3.095 0.925 ;
        RECT 3.785 0.755 3.955 0.925 ;
        RECT 4.645 0.755 4.815 0.925 ;
        RECT 7.225 0.755 7.395 0.925 ;
        RECT 8.085 0.755 8.255 0.925 ;
        RECT 8.945 0.755 9.115 0.925 ;
        RECT 9.805 0.755 9.975 0.925 ;
        RECT 10.665 0.755 10.835 0.925 ;
      LAYER met1 ;
        RECT 4.130 29.260 7.910 29.540 ;
        RECT 4.130 27.160 7.910 27.440 ;
        RECT 3.700 23.380 8.340 23.660 ;
        RECT 4.130 22.960 7.910 23.240 ;
        RECT 3.280 22.540 5.750 22.820 ;
        RECT 4.130 22.120 7.910 22.400 ;
        RECT 3.700 21.700 8.340 21.980 ;
        RECT 5.430 21.280 8.330 21.560 ;
        RECT 4.130 17.920 7.910 18.200 ;
        RECT 4.130 15.820 7.910 16.100 ;
        RECT 1.120 14.140 4.900 14.420 ;
        RECT 7.140 14.140 10.920 14.420 ;
        RECT 1.120 12.040 4.900 12.320 ;
        RECT 7.140 12.040 10.920 12.320 ;
        RECT 3.280 11.200 8.760 11.480 ;
        RECT 0.690 8.260 5.330 8.540 ;
        RECT 6.710 8.260 11.350 8.540 ;
        RECT 1.120 7.840 4.900 8.120 ;
        RECT 7.140 7.840 10.920 8.120 ;
        RECT 4.570 7.420 6.190 7.700 ;
        RECT 8.010 7.420 8.760 7.700 ;
        RECT 1.120 7.000 4.900 7.280 ;
        RECT 5.850 7.000 10.920 7.280 ;
        RECT 0.690 6.580 5.330 6.860 ;
        RECT 6.710 6.580 11.350 6.860 ;
        RECT 3.280 3.640 8.760 3.920 ;
        RECT 1.120 2.800 4.900 3.080 ;
        RECT 7.140 2.800 10.920 3.080 ;
        RECT 1.120 0.700 4.900 0.980 ;
        RECT 7.140 0.700 10.920 0.980 ;
      LAYER via ;
        RECT 5.460 29.270 5.720 29.530 ;
        RECT 6.320 27.170 6.580 27.430 ;
        RECT 5.460 23.390 5.720 23.650 ;
        RECT 5.890 22.970 6.150 23.230 ;
        RECT 3.310 22.550 3.570 22.810 ;
        RECT 5.460 22.550 5.720 22.810 ;
        RECT 5.890 22.130 6.150 22.390 ;
        RECT 7.180 22.130 7.440 22.390 ;
        RECT 5.460 21.710 5.720 21.970 ;
        RECT 5.460 21.290 5.720 21.550 ;
        RECT 8.040 21.290 8.300 21.550 ;
        RECT 4.170 17.930 4.430 18.190 ;
        RECT 6.320 17.930 6.580 18.190 ;
        RECT 5.460 15.830 5.720 16.090 ;
        RECT 3.310 14.150 3.570 14.410 ;
        RECT 8.470 14.150 8.730 14.410 ;
        RECT 4.600 12.050 4.860 12.310 ;
        RECT 7.180 12.050 7.440 12.310 ;
        RECT 8.900 12.050 9.160 12.310 ;
        RECT 3.310 11.210 3.570 11.470 ;
        RECT 8.470 11.210 8.730 11.470 ;
        RECT 3.310 8.270 3.570 8.530 ;
        RECT 8.470 8.270 8.730 8.530 ;
        RECT 2.880 7.850 3.140 8.110 ;
        RECT 4.170 7.850 4.430 8.110 ;
        RECT 7.180 7.850 7.440 8.110 ;
        RECT 4.600 7.430 4.860 7.690 ;
        RECT 8.040 7.430 8.300 7.690 ;
        RECT 8.470 7.430 8.730 7.690 ;
        RECT 2.880 7.010 3.140 7.270 ;
        RECT 7.180 7.010 7.440 7.270 ;
        RECT 3.310 6.590 3.570 6.850 ;
        RECT 8.470 6.590 8.730 6.850 ;
        RECT 3.310 3.650 3.570 3.910 ;
        RECT 8.470 3.650 8.730 3.910 ;
        RECT 4.600 2.810 4.860 3.070 ;
        RECT 8.900 2.810 9.160 3.070 ;
        RECT 3.310 0.710 3.570 0.970 ;
        RECT 8.470 0.710 8.730 0.970 ;
      LAYER met2 ;
        RECT 3.300 8.240 3.580 22.840 ;
        RECT 5.450 22.520 5.730 29.560 ;
        RECT 5.880 22.100 6.160 23.260 ;
        RECT 2.870 6.980 3.150 8.140 ;
        RECT 4.160 7.820 4.440 18.220 ;
        RECT 5.450 15.800 5.730 22.000 ;
        RECT 6.310 17.900 6.590 27.460 ;
        RECT 3.300 0.680 3.580 6.880 ;
        RECT 4.590 2.780 4.870 12.340 ;
        RECT 7.170 12.020 7.450 22.420 ;
        RECT 7.170 6.980 7.450 8.140 ;
        RECT 8.030 7.400 8.310 21.580 ;
        RECT 8.460 8.240 8.740 14.440 ;
        RECT 8.460 0.680 8.740 7.720 ;
        RECT 8.890 2.780 9.170 12.340 ;
  END
END RINGOSC_0
END LIBRARY

