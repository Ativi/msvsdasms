module RingOsc_cap (
        output out
);


endmodule
