module adc (
      input vin,
      input vref,
      output out
);


endmodule
