MACRO ONEBITADC
  ORIGIN 0 0 ;
  FOREIGN ONEBITADC 0 0 ;
  SIZE 15.48 BY 22.68 ;
  PIN OUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 8.86 15.82 13.5 16.1 ;
      LAYER M2 ;
        RECT 11.44 14.56 14.36 14.84 ;
      LAYER M2 ;
        RECT 11.88 15.82 12.2 16.1 ;
      LAYER M3 ;
        RECT 11.9 14.7 12.18 15.96 ;
      LAYER M2 ;
        RECT 11.88 14.56 12.2 14.84 ;
    END
  END OUT
  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 9.75 0.68 10.03 6.46 ;
      LAYER M3 ;
        RECT 8.03 8.24 8.31 14.44 ;
      LAYER M3 ;
        RECT 12.33 8.24 12.61 14.44 ;
      LAYER M3 ;
        RECT 9.75 6.3 10.03 7.98 ;
      LAYER M2 ;
        RECT 8.17 7.84 9.89 8.12 ;
      LAYER M3 ;
        RECT 8.03 7.98 8.31 8.4 ;
      LAYER M2 ;
        RECT 9.89 7.84 12.47 8.12 ;
      LAYER M3 ;
        RECT 12.33 7.98 12.61 8.4 ;
    END
  END VDD
  PIN VIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.12 12.04 4.04 12.32 ;
    END
  END VIN
  PIN VREF
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.12 2.8 4.04 3.08 ;
    END
  END VREF
  OBS 
  LAYER M3 ;
        RECT 7.6 10.34 7.88 14.86 ;
  LAYER M2 ;
        RECT 2.84 19.6 5.76 19.88 ;
  LAYER M3 ;
        RECT 10.61 15.38 10.89 19.9 ;
  LAYER M2 ;
        RECT 5.59 19.6 7.31 19.88 ;
  LAYER M3 ;
        RECT 7.17 19.32 7.45 19.74 ;
  LAYER M2 ;
        RECT 7.31 19.18 10.75 19.46 ;
  LAYER M3 ;
        RECT 10.61 19.135 10.89 19.505 ;
  LAYER M3 ;
        RECT 7.6 14.7 7.88 15.12 ;
  LAYER M2 ;
        RECT 7.74 14.98 10.75 15.26 ;
  LAYER M3 ;
        RECT 10.61 15.12 10.89 15.54 ;
  LAYER M2 ;
        RECT 7.58 14.98 7.9 15.26 ;
  LAYER M3 ;
        RECT 7.6 14.96 7.88 15.28 ;
  LAYER M2 ;
        RECT 10.59 14.98 10.91 15.26 ;
  LAYER M3 ;
        RECT 10.61 14.96 10.89 15.28 ;
  LAYER M2 ;
        RECT 7.58 14.98 7.9 15.26 ;
  LAYER M3 ;
        RECT 7.6 14.96 7.88 15.28 ;
  LAYER M2 ;
        RECT 10.59 14.98 10.91 15.26 ;
  LAYER M3 ;
        RECT 10.61 14.96 10.89 15.28 ;
  LAYER M3 ;
        RECT 2.87 0.68 3.15 6.88 ;
  LAYER M3 ;
        RECT 2.87 8.24 3.15 14.44 ;
  LAYER M2 ;
        RECT 2.84 15.4 5.76 15.68 ;
  LAYER M3 ;
        RECT 2.87 6.72 3.15 8.4 ;
  LAYER M3 ;
        RECT 2.87 14.28 3.15 15.54 ;
  LAYER M2 ;
        RECT 2.85 15.4 3.17 15.68 ;
  LAYER M2 ;
        RECT 2.85 15.4 3.17 15.68 ;
  LAYER M3 ;
        RECT 2.87 15.38 3.15 15.7 ;
  LAYER M2 ;
        RECT 2.85 15.4 3.17 15.68 ;
  LAYER M3 ;
        RECT 2.87 15.38 3.15 15.7 ;
  LAYER M3 ;
        RECT 4.59 15.8 4.87 22 ;
  LAYER M3 ;
        RECT 11.47 16.22 11.75 22 ;
  LAYER M3 ;
        RECT 4.59 18.715 4.87 19.085 ;
  LAYER M2 ;
        RECT 4.73 18.76 11.61 19.04 ;
  LAYER M3 ;
        RECT 11.47 18.715 11.75 19.085 ;
  LAYER M2 ;
        RECT 1.12 7 4.04 7.28 ;
  LAYER M3 ;
        RECT 8.89 2.78 9.17 7.3 ;
  LAYER M2 ;
        RECT 3.87 7 5.59 7.28 ;
  LAYER M3 ;
        RECT 5.45 6.3 5.73 7.14 ;
  LAYER M4 ;
        RECT 5.59 5.9 9.03 6.7 ;
  LAYER M3 ;
        RECT 8.89 6.115 9.17 6.485 ;
  LAYER M2 ;
        RECT 5.43 7 5.75 7.28 ;
  LAYER M3 ;
        RECT 5.45 6.98 5.73 7.3 ;
  LAYER M3 ;
        RECT 5.45 6.115 5.73 6.485 ;
  LAYER M4 ;
        RECT 5.425 5.9 5.755 6.7 ;
  LAYER M3 ;
        RECT 8.89 6.115 9.17 6.485 ;
  LAYER M4 ;
        RECT 8.865 5.9 9.195 6.7 ;
  LAYER M2 ;
        RECT 5.43 7 5.75 7.28 ;
  LAYER M3 ;
        RECT 5.45 6.98 5.73 7.3 ;
  LAYER M3 ;
        RECT 5.45 6.115 5.73 6.485 ;
  LAYER M4 ;
        RECT 5.425 5.9 5.755 6.7 ;
  LAYER M3 ;
        RECT 8.89 6.115 9.17 6.485 ;
  LAYER M4 ;
        RECT 8.865 5.9 9.195 6.7 ;
  LAYER M2 ;
        RECT 1.12 7.84 4.04 8.12 ;
  LAYER M2 ;
        RECT 7.14 6.58 11.78 6.86 ;
  LAYER M2 ;
        RECT 11.44 10.36 14.36 10.64 ;
  LAYER M2 ;
        RECT 3.87 7.84 7.31 8.12 ;
  LAYER M3 ;
        RECT 7.17 6.72 7.45 7.98 ;
  LAYER M2 ;
        RECT 7.15 6.58 7.47 6.86 ;
  LAYER M2 ;
        RECT 11.45 6.58 11.77 6.86 ;
  LAYER M3 ;
        RECT 11.47 6.72 11.75 10.5 ;
  LAYER M2 ;
        RECT 11.45 10.36 11.77 10.64 ;
  LAYER M2 ;
        RECT 7.15 6.58 7.47 6.86 ;
  LAYER M3 ;
        RECT 7.17 6.56 7.45 6.88 ;
  LAYER M2 ;
        RECT 7.15 7.84 7.47 8.12 ;
  LAYER M3 ;
        RECT 7.17 7.82 7.45 8.14 ;
  LAYER M2 ;
        RECT 7.15 6.58 7.47 6.86 ;
  LAYER M3 ;
        RECT 7.17 6.56 7.45 6.88 ;
  LAYER M2 ;
        RECT 7.15 7.84 7.47 8.12 ;
  LAYER M3 ;
        RECT 7.17 7.82 7.45 8.14 ;
  LAYER M2 ;
        RECT 7.15 6.58 7.47 6.86 ;
  LAYER M3 ;
        RECT 7.17 6.56 7.45 6.88 ;
  LAYER M2 ;
        RECT 7.15 7.84 7.47 8.12 ;
  LAYER M3 ;
        RECT 7.17 7.82 7.45 8.14 ;
  LAYER M2 ;
        RECT 11.45 6.58 11.77 6.86 ;
  LAYER M3 ;
        RECT 11.47 6.56 11.75 6.88 ;
  LAYER M2 ;
        RECT 11.45 10.36 11.77 10.64 ;
  LAYER M3 ;
        RECT 11.47 10.34 11.75 10.66 ;
  LAYER M2 ;
        RECT 7.15 6.58 7.47 6.86 ;
  LAYER M3 ;
        RECT 7.17 6.56 7.45 6.88 ;
  LAYER M2 ;
        RECT 7.15 7.84 7.47 8.12 ;
  LAYER M3 ;
        RECT 7.17 7.82 7.45 8.14 ;
  LAYER M2 ;
        RECT 11.45 6.58 11.77 6.86 ;
  LAYER M3 ;
        RECT 11.47 6.56 11.75 6.88 ;
  LAYER M2 ;
        RECT 11.45 10.36 11.77 10.64 ;
  LAYER M3 ;
        RECT 11.47 10.34 11.75 10.66 ;
  LAYER M1 ;
        RECT 8.045 15.455 8.295 18.985 ;
  LAYER M1 ;
        RECT 8.045 19.235 8.295 20.245 ;
  LAYER M1 ;
        RECT 8.045 21.335 8.295 22.345 ;
  LAYER M1 ;
        RECT 7.615 15.455 7.865 18.985 ;
  LAYER M1 ;
        RECT 8.475 15.455 8.725 18.985 ;
  LAYER M1 ;
        RECT 8.905 15.455 9.155 18.985 ;
  LAYER M1 ;
        RECT 8.905 19.235 9.155 20.245 ;
  LAYER M1 ;
        RECT 8.905 21.335 9.155 22.345 ;
  LAYER M1 ;
        RECT 9.335 15.455 9.585 18.985 ;
  LAYER M1 ;
        RECT 9.765 15.455 10.015 18.985 ;
  LAYER M1 ;
        RECT 9.765 19.235 10.015 20.245 ;
  LAYER M1 ;
        RECT 9.765 21.335 10.015 22.345 ;
  LAYER M1 ;
        RECT 10.195 15.455 10.445 18.985 ;
  LAYER M1 ;
        RECT 10.625 15.455 10.875 18.985 ;
  LAYER M1 ;
        RECT 10.625 19.235 10.875 20.245 ;
  LAYER M1 ;
        RECT 10.625 21.335 10.875 22.345 ;
  LAYER M1 ;
        RECT 11.055 15.455 11.305 18.985 ;
  LAYER M1 ;
        RECT 11.485 15.455 11.735 18.985 ;
  LAYER M1 ;
        RECT 11.485 19.235 11.735 20.245 ;
  LAYER M1 ;
        RECT 11.485 21.335 11.735 22.345 ;
  LAYER M1 ;
        RECT 11.915 15.455 12.165 18.985 ;
  LAYER M1 ;
        RECT 12.345 15.455 12.595 18.985 ;
  LAYER M1 ;
        RECT 12.345 19.235 12.595 20.245 ;
  LAYER M1 ;
        RECT 12.345 21.335 12.595 22.345 ;
  LAYER M1 ;
        RECT 12.775 15.455 13.025 18.985 ;
  LAYER M1 ;
        RECT 13.205 15.455 13.455 18.985 ;
  LAYER M1 ;
        RECT 13.205 19.235 13.455 20.245 ;
  LAYER M1 ;
        RECT 13.205 21.335 13.455 22.345 ;
  LAYER M1 ;
        RECT 13.635 15.455 13.885 18.985 ;
  LAYER M1 ;
        RECT 14.065 15.455 14.315 18.985 ;
  LAYER M1 ;
        RECT 14.065 19.235 14.315 20.245 ;
  LAYER M1 ;
        RECT 14.065 21.335 14.315 22.345 ;
  LAYER M1 ;
        RECT 14.495 15.455 14.745 18.985 ;
  LAYER M2 ;
        RECT 8 19.6 14.36 19.88 ;
  LAYER M2 ;
        RECT 8 15.4 14.36 15.68 ;
  LAYER M2 ;
        RECT 8 21.7 14.36 21.98 ;
  LAYER M2 ;
        RECT 7.57 16.24 14.79 16.52 ;
  LAYER M3 ;
        RECT 10.61 15.38 10.89 19.9 ;
  LAYER M2 ;
        RECT 8.86 15.82 13.5 16.1 ;
  LAYER M3 ;
        RECT 11.47 16.22 11.75 22 ;
  LAYER M1 ;
        RECT 2.885 15.455 3.135 18.985 ;
  LAYER M1 ;
        RECT 2.885 19.235 3.135 20.245 ;
  LAYER M1 ;
        RECT 2.885 21.335 3.135 22.345 ;
  LAYER M1 ;
        RECT 2.455 15.455 2.705 18.985 ;
  LAYER M1 ;
        RECT 3.315 15.455 3.565 18.985 ;
  LAYER M1 ;
        RECT 3.745 15.455 3.995 18.985 ;
  LAYER M1 ;
        RECT 3.745 19.235 3.995 20.245 ;
  LAYER M1 ;
        RECT 3.745 21.335 3.995 22.345 ;
  LAYER M1 ;
        RECT 4.175 15.455 4.425 18.985 ;
  LAYER M1 ;
        RECT 4.605 15.455 4.855 18.985 ;
  LAYER M1 ;
        RECT 4.605 19.235 4.855 20.245 ;
  LAYER M1 ;
        RECT 4.605 21.335 4.855 22.345 ;
  LAYER M1 ;
        RECT 5.035 15.455 5.285 18.985 ;
  LAYER M1 ;
        RECT 5.465 15.455 5.715 18.985 ;
  LAYER M1 ;
        RECT 5.465 19.235 5.715 20.245 ;
  LAYER M1 ;
        RECT 5.465 21.335 5.715 22.345 ;
  LAYER M1 ;
        RECT 5.895 15.455 6.145 18.985 ;
  LAYER M2 ;
        RECT 2.84 21.7 5.76 21.98 ;
  LAYER M2 ;
        RECT 2.41 15.82 6.19 16.1 ;
  LAYER M2 ;
        RECT 2.84 15.4 5.76 15.68 ;
  LAYER M2 ;
        RECT 2.84 19.6 5.76 19.88 ;
  LAYER M3 ;
        RECT 4.59 15.8 4.87 22 ;
  LAYER M1 ;
        RECT 6.325 3.695 6.575 7.225 ;
  LAYER M1 ;
        RECT 6.325 2.435 6.575 3.445 ;
  LAYER M1 ;
        RECT 6.325 0.335 6.575 1.345 ;
  LAYER M1 ;
        RECT 5.895 3.695 6.145 7.225 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M1 ;
        RECT 7.185 3.695 7.435 7.225 ;
  LAYER M1 ;
        RECT 7.185 2.435 7.435 3.445 ;
  LAYER M1 ;
        RECT 7.185 0.335 7.435 1.345 ;
  LAYER M1 ;
        RECT 7.615 3.695 7.865 7.225 ;
  LAYER M1 ;
        RECT 8.045 3.695 8.295 7.225 ;
  LAYER M1 ;
        RECT 8.045 2.435 8.295 3.445 ;
  LAYER M1 ;
        RECT 8.045 0.335 8.295 1.345 ;
  LAYER M1 ;
        RECT 8.475 3.695 8.725 7.225 ;
  LAYER M1 ;
        RECT 8.905 3.695 9.155 7.225 ;
  LAYER M1 ;
        RECT 8.905 2.435 9.155 3.445 ;
  LAYER M1 ;
        RECT 8.905 0.335 9.155 1.345 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M1 ;
        RECT 9.765 3.695 10.015 7.225 ;
  LAYER M1 ;
        RECT 9.765 2.435 10.015 3.445 ;
  LAYER M1 ;
        RECT 9.765 0.335 10.015 1.345 ;
  LAYER M1 ;
        RECT 10.195 3.695 10.445 7.225 ;
  LAYER M1 ;
        RECT 10.625 3.695 10.875 7.225 ;
  LAYER M1 ;
        RECT 10.625 2.435 10.875 3.445 ;
  LAYER M1 ;
        RECT 10.625 0.335 10.875 1.345 ;
  LAYER M1 ;
        RECT 11.055 3.695 11.305 7.225 ;
  LAYER M1 ;
        RECT 11.485 3.695 11.735 7.225 ;
  LAYER M1 ;
        RECT 11.485 2.435 11.735 3.445 ;
  LAYER M1 ;
        RECT 11.485 0.335 11.735 1.345 ;
  LAYER M1 ;
        RECT 11.915 3.695 12.165 7.225 ;
  LAYER M1 ;
        RECT 12.345 3.695 12.595 7.225 ;
  LAYER M1 ;
        RECT 12.345 2.435 12.595 3.445 ;
  LAYER M1 ;
        RECT 12.345 0.335 12.595 1.345 ;
  LAYER M1 ;
        RECT 12.775 3.695 13.025 7.225 ;
  LAYER M2 ;
        RECT 6.28 2.8 12.64 3.08 ;
  LAYER M2 ;
        RECT 6.28 7 12.64 7.28 ;
  LAYER M2 ;
        RECT 6.28 0.7 12.64 0.98 ;
  LAYER M2 ;
        RECT 5.85 6.16 13.07 6.44 ;
  LAYER M3 ;
        RECT 8.89 2.78 9.17 7.3 ;
  LAYER M2 ;
        RECT 7.14 6.58 11.78 6.86 ;
  LAYER M3 ;
        RECT 9.75 0.68 10.03 6.46 ;
  LAYER M1 ;
        RECT 6.325 11.255 6.575 14.785 ;
  LAYER M1 ;
        RECT 6.325 9.995 6.575 11.005 ;
  LAYER M1 ;
        RECT 6.325 7.895 6.575 8.905 ;
  LAYER M1 ;
        RECT 5.895 11.255 6.145 14.785 ;
  LAYER M1 ;
        RECT 6.755 11.255 7.005 14.785 ;
  LAYER M1 ;
        RECT 7.185 11.255 7.435 14.785 ;
  LAYER M1 ;
        RECT 7.185 9.995 7.435 11.005 ;
  LAYER M1 ;
        RECT 7.185 7.895 7.435 8.905 ;
  LAYER M1 ;
        RECT 7.615 11.255 7.865 14.785 ;
  LAYER M1 ;
        RECT 8.045 11.255 8.295 14.785 ;
  LAYER M1 ;
        RECT 8.045 9.995 8.295 11.005 ;
  LAYER M1 ;
        RECT 8.045 7.895 8.295 8.905 ;
  LAYER M1 ;
        RECT 8.475 11.255 8.725 14.785 ;
  LAYER M1 ;
        RECT 8.905 11.255 9.155 14.785 ;
  LAYER M1 ;
        RECT 8.905 9.995 9.155 11.005 ;
  LAYER M1 ;
        RECT 8.905 7.895 9.155 8.905 ;
  LAYER M1 ;
        RECT 9.335 11.255 9.585 14.785 ;
  LAYER M2 ;
        RECT 6.28 10.36 9.2 10.64 ;
  LAYER M2 ;
        RECT 6.28 14.56 9.2 14.84 ;
  LAYER M2 ;
        RECT 6.28 8.26 9.2 8.54 ;
  LAYER M2 ;
        RECT 5.85 14.14 9.63 14.42 ;
  LAYER M3 ;
        RECT 7.6 10.34 7.88 14.86 ;
  LAYER M3 ;
        RECT 8.03 8.24 8.31 14.44 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 11.425 ;
  LAYER M1 ;
        RECT 1.165 11.675 1.415 12.685 ;
  LAYER M1 ;
        RECT 1.165 13.775 1.415 14.785 ;
  LAYER M1 ;
        RECT 0.735 7.895 0.985 11.425 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 11.425 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 11.425 ;
  LAYER M1 ;
        RECT 2.025 11.675 2.275 12.685 ;
  LAYER M1 ;
        RECT 2.025 13.775 2.275 14.785 ;
  LAYER M1 ;
        RECT 2.455 7.895 2.705 11.425 ;
  LAYER M1 ;
        RECT 2.885 7.895 3.135 11.425 ;
  LAYER M1 ;
        RECT 2.885 11.675 3.135 12.685 ;
  LAYER M1 ;
        RECT 2.885 13.775 3.135 14.785 ;
  LAYER M1 ;
        RECT 3.315 7.895 3.565 11.425 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 11.425 ;
  LAYER M1 ;
        RECT 3.745 11.675 3.995 12.685 ;
  LAYER M1 ;
        RECT 3.745 13.775 3.995 14.785 ;
  LAYER M1 ;
        RECT 4.175 7.895 4.425 11.425 ;
  LAYER M2 ;
        RECT 1.12 14.14 4.04 14.42 ;
  LAYER M2 ;
        RECT 0.69 8.26 4.47 8.54 ;
  LAYER M2 ;
        RECT 1.12 7.84 4.04 8.12 ;
  LAYER M2 ;
        RECT 1.12 12.04 4.04 12.32 ;
  LAYER M3 ;
        RECT 2.87 8.24 3.15 14.44 ;
  LAYER M1 ;
        RECT 1.165 3.695 1.415 7.225 ;
  LAYER M1 ;
        RECT 1.165 2.435 1.415 3.445 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 1.345 ;
  LAYER M1 ;
        RECT 0.735 3.695 0.985 7.225 ;
  LAYER M1 ;
        RECT 1.595 3.695 1.845 7.225 ;
  LAYER M1 ;
        RECT 2.025 3.695 2.275 7.225 ;
  LAYER M1 ;
        RECT 2.025 2.435 2.275 3.445 ;
  LAYER M1 ;
        RECT 2.025 0.335 2.275 1.345 ;
  LAYER M1 ;
        RECT 2.455 3.695 2.705 7.225 ;
  LAYER M1 ;
        RECT 2.885 3.695 3.135 7.225 ;
  LAYER M1 ;
        RECT 2.885 2.435 3.135 3.445 ;
  LAYER M1 ;
        RECT 2.885 0.335 3.135 1.345 ;
  LAYER M1 ;
        RECT 3.315 3.695 3.565 7.225 ;
  LAYER M1 ;
        RECT 3.745 3.695 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.745 2.435 3.995 3.445 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 1.345 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M2 ;
        RECT 1.12 0.7 4.04 0.98 ;
  LAYER M2 ;
        RECT 0.69 6.58 4.47 6.86 ;
  LAYER M2 ;
        RECT 1.12 7 4.04 7.28 ;
  LAYER M2 ;
        RECT 1.12 2.8 4.04 3.08 ;
  LAYER M3 ;
        RECT 2.87 0.68 3.15 6.88 ;
  LAYER M1 ;
        RECT 14.065 11.255 14.315 14.785 ;
  LAYER M1 ;
        RECT 14.065 9.995 14.315 11.005 ;
  LAYER M1 ;
        RECT 14.065 7.895 14.315 8.905 ;
  LAYER M1 ;
        RECT 14.495 11.255 14.745 14.785 ;
  LAYER M1 ;
        RECT 13.635 11.255 13.885 14.785 ;
  LAYER M1 ;
        RECT 13.205 11.255 13.455 14.785 ;
  LAYER M1 ;
        RECT 13.205 9.995 13.455 11.005 ;
  LAYER M1 ;
        RECT 13.205 7.895 13.455 8.905 ;
  LAYER M1 ;
        RECT 12.775 11.255 13.025 14.785 ;
  LAYER M1 ;
        RECT 12.345 11.255 12.595 14.785 ;
  LAYER M1 ;
        RECT 12.345 9.995 12.595 11.005 ;
  LAYER M1 ;
        RECT 12.345 7.895 12.595 8.905 ;
  LAYER M1 ;
        RECT 11.915 11.255 12.165 14.785 ;
  LAYER M1 ;
        RECT 11.485 11.255 11.735 14.785 ;
  LAYER M1 ;
        RECT 11.485 9.995 11.735 11.005 ;
  LAYER M1 ;
        RECT 11.485 7.895 11.735 8.905 ;
  LAYER M1 ;
        RECT 11.055 11.255 11.305 14.785 ;
  LAYER M2 ;
        RECT 11.44 8.26 14.36 8.54 ;
  LAYER M2 ;
        RECT 11.01 14.14 14.79 14.42 ;
  LAYER M2 ;
        RECT 11.44 14.56 14.36 14.84 ;
  LAYER M2 ;
        RECT 11.44 10.36 14.36 10.64 ;
  LAYER M3 ;
        RECT 12.33 8.24 12.61 14.44 ;
  END 
END ONEBITADC
