module analog_async_up_down (Vin,
    out,
    vref);
 output Vin;
 output out;
 input vref;


 sky130_fd_sc_hd__conb_1 _1_ (.LO(Vin));
 sky130_fd_sc_hd__conb_1 _3_ (.LO(out));
 sky130_fd_sc_hd__decap_4 PHY_0 ();
 sky130_fd_sc_hd__decap_4 PHY_1 ();
 sky130_fd_sc_hd__decap_4 PHY_2 ();
 sky130_fd_sc_hd__decap_4 PHY_3 ();
 sky130_fd_sc_hd__decap_4 PHY_4 ();
 sky130_fd_sc_hd__decap_4 PHY_5 ();
 sky130_fd_sc_hd__decap_4 PHY_6 ();
 sky130_fd_sc_hd__decap_4 PHY_7 ();
 sky130_fd_sc_hd__decap_4 PHY_8 ();
 sky130_fd_sc_hd__decap_4 PHY_9 ();
 sky130_fd_sc_hd__decap_4 PHY_10 ();
 sky130_fd_sc_hd__decap_4 PHY_11 ();
 sky130_fd_sc_hd__decap_4 PHY_12 ();
 sky130_fd_sc_hd__decap_4 PHY_13 ();
 sky130_fd_sc_hd__decap_4 PHY_14 ();
 sky130_fd_sc_hd__decap_4 PHY_15 ();
 sky130_fd_sc_hd__decap_4 PHY_16 ();
 sky130_fd_sc_hd__decap_4 PHY_17 ();
 sky130_fd_sc_hd__decap_4 PHY_18 ();
 sky130_fd_sc_hd__decap_4 PHY_19 ();
 sky130_fd_sc_hd__decap_4 PHY_20 ();
 sky130_fd_sc_hd__decap_4 PHY_21 ();
 sky130_fd_sc_hd__decap_4 PHY_22 ();
 sky130_fd_sc_hd__decap_4 PHY_23 ();
 sky130_fd_sc_hd__decap_4 PHY_24 ();
 sky130_fd_sc_hd__decap_4 PHY_25 ();
 sky130_fd_sc_hd__decap_4 PHY_26 ();
 sky130_fd_sc_hd__decap_4 PHY_27 ();
 sky130_fd_sc_hd__decap_4 PHY_28 ();
 sky130_fd_sc_hd__decap_4 PHY_29 ();
 sky130_fd_sc_hd__decap_4 PHY_30 ();
 sky130_fd_sc_hd__decap_4 PHY_31 ();
 sky130_fd_sc_hd__decap_4 PHY_32 ();
 sky130_fd_sc_hd__decap_4 PHY_33 ();
 sky130_fd_sc_hd__decap_4 PHY_34 ();
 sky130_fd_sc_hd__decap_4 PHY_35 ();
 sky130_fd_sc_hd__decap_4 PHY_36 ();
 sky130_fd_sc_hd__decap_4 PHY_37 ();
 sky130_fd_sc_hd__decap_4 PHY_38 ();
 sky130_fd_sc_hd__decap_4 PHY_39 ();
 sky130_fd_sc_hd__decap_4 PHY_40 ();
 sky130_fd_sc_hd__decap_4 PHY_41 ();
 sky130_fd_sc_hd__decap_4 PHY_42 ();
 sky130_fd_sc_hd__decap_4 PHY_43 ();
 sky130_fd_sc_hd__decap_4 PHY_44 ();
 sky130_fd_sc_hd__decap_4 PHY_45 ();
 sky130_fd_sc_hd__decap_4 PHY_46 ();
 sky130_fd_sc_hd__decap_4 PHY_47 ();
 sky130_fd_sc_hd__decap_4 PHY_48 ();
 sky130_fd_sc_hd__decap_4 PHY_49 ();
 sky130_fd_sc_hd__decap_4 PHY_50 ();
 sky130_fd_sc_hd__decap_4 PHY_51 ();
 sky130_fd_sc_hd__decap_4 PHY_52 ();
 sky130_fd_sc_hd__decap_4 PHY_53 ();
 sky130_fd_sc_hd__decap_4 PHY_54 ();
 sky130_fd_sc_hd__decap_4 PHY_55 ();
 sky130_fd_sc_hd__decap_4 PHY_56 ();
 sky130_fd_sc_hd__decap_4 PHY_57 ();
 sky130_fd_sc_hd__decap_4 PHY_58 ();
 sky130_fd_sc_hd__decap_4 PHY_59 ();
 sky130_fd_sc_hd__decap_4 PHY_60 ();
 sky130_fd_sc_hd__decap_4 PHY_61 ();
 sky130_fd_sc_hd__decap_4 PHY_62 ();
 sky130_fd_sc_hd__decap_4 PHY_63 ();
 sky130_fd_sc_hd__decap_4 PHY_64 ();
 sky130_fd_sc_hd__decap_4 PHY_65 ();
 sky130_fd_sc_hd__decap_4 PHY_66 ();
 sky130_fd_sc_hd__decap_4 PHY_67 ();
 sky130_fd_sc_hd__decap_4 PHY_68 ();
 sky130_fd_sc_hd__decap_4 PHY_69 ();
 sky130_fd_sc_hd__decap_4 PHY_70 ();
 sky130_fd_sc_hd__decap_4 PHY_71 ();
 sky130_fd_sc_hd__decap_4 PHY_72 ();
 sky130_fd_sc_hd__decap_4 PHY_73 ();
 sky130_fd_sc_hd__decap_4 PHY_74 ();
 sky130_fd_sc_hd__decap_4 PHY_75 ();
 sky130_fd_sc_hd__decap_4 PHY_76 ();
 sky130_fd_sc_hd__decap_4 PHY_77 ();
 sky130_fd_sc_hd__decap_4 PHY_78 ();
 sky130_fd_sc_hd__decap_4 PHY_79 ();
 sky130_fd_sc_hd__decap_4 PHY_80 ();
 sky130_fd_sc_hd__decap_4 PHY_81 ();
 sky130_fd_sc_hd__decap_4 PHY_82 ();
 sky130_fd_sc_hd__decap_4 PHY_83 ();
 sky130_fd_sc_hd__decap_4 PHY_84 ();
 sky130_fd_sc_hd__decap_4 PHY_85 ();
 sky130_fd_sc_hd__decap_4 PHY_86 ();
 sky130_fd_sc_hd__decap_4 PHY_87 ();
 sky130_fd_sc_hd__decap_4 PHY_88 ();
 sky130_fd_sc_hd__decap_4 PHY_89 ();
 sky130_fd_sc_hd__decap_4 PHY_90 ();
 sky130_fd_sc_hd__decap_4 PHY_91 ();
 sky130_fd_sc_hd__decap_4 PHY_92 ();
 sky130_fd_sc_hd__decap_4 PHY_93 ();
 sky130_fd_sc_hd__decap_4 PHY_94 ();
 sky130_fd_sc_hd__decap_4 PHY_95 ();
 sky130_fd_sc_hd__decap_4 PHY_96 ();
 sky130_fd_sc_hd__decap_4 PHY_97 ();
 sky130_fd_sc_hd__decap_4 PHY_98 ();
 sky130_fd_sc_hd__decap_4 PHY_99 ();
 sky130_fd_sc_hd__decap_4 PHY_100 ();
 sky130_fd_sc_hd__decap_4 PHY_101 ();
 sky130_fd_sc_hd__decap_4 PHY_102 ();
 sky130_fd_sc_hd__decap_4 PHY_103 ();
 sky130_fd_sc_hd__decap_4 PHY_104 ();
 sky130_fd_sc_hd__decap_4 PHY_105 ();
 sky130_fd_sc_hd__decap_4 PHY_106 ();
 sky130_fd_sc_hd__decap_4 PHY_107 ();
 sky130_fd_sc_hd__decap_4 PHY_108 ();
 sky130_fd_sc_hd__decap_4 PHY_109 ();
 sky130_fd_sc_hd__decap_4 PHY_110 ();
 sky130_fd_sc_hd__decap_4 PHY_111 ();
 sky130_fd_sc_hd__decap_4 PHY_112 ();
 sky130_fd_sc_hd__decap_4 PHY_113 ();
 sky130_fd_sc_hd__decap_4 PHY_114 ();
 sky130_fd_sc_hd__decap_4 PHY_115 ();
 sky130_fd_sc_hd__decap_4 PHY_116 ();
 sky130_fd_sc_hd__decap_4 PHY_117 ();
 sky130_fd_sc_hd__decap_4 PHY_118 ();
 sky130_fd_sc_hd__decap_4 PHY_119 ();
 sky130_fd_sc_hd__decap_4 PHY_120 ();
 sky130_fd_sc_hd__decap_4 PHY_121 ();
 sky130_fd_sc_hd__decap_4 PHY_122 ();
 sky130_fd_sc_hd__decap_4 PHY_123 ();
 sky130_fd_sc_hd__decap_4 PHY_124 ();
 sky130_fd_sc_hd__decap_4 PHY_125 ();
 sky130_fd_sc_hd__decap_4 PHY_126 ();
 sky130_fd_sc_hd__decap_4 PHY_127 ();
 sky130_fd_sc_hd__decap_4 PHY_128 ();
 sky130_fd_sc_hd__decap_4 PHY_129 ();
 sky130_fd_sc_hd__decap_4 PHY_130 ();
 sky130_fd_sc_hd__decap_4 PHY_131 ();
 sky130_fd_sc_hd__decap_4 PHY_132 ();
 sky130_fd_sc_hd__decap_4 PHY_133 ();
 sky130_fd_sc_hd__decap_4 PHY_134 ();
 sky130_fd_sc_hd__decap_4 PHY_135 ();
 sky130_fd_sc_hd__decap_4 PHY_136 ();
 sky130_fd_sc_hd__decap_4 PHY_137 ();
 sky130_fd_sc_hd__decap_4 PHY_138 ();
 sky130_fd_sc_hd__decap_4 PHY_139 ();
 sky130_fd_sc_hd__decap_4 PHY_140 ();
 sky130_fd_sc_hd__decap_4 PHY_141 ();
 sky130_fd_sc_hd__decap_4 PHY_142 ();
 sky130_fd_sc_hd__decap_4 PHY_143 ();
 sky130_fd_sc_hd__decap_4 PHY_144 ();
 sky130_fd_sc_hd__decap_4 PHY_145 ();
 sky130_fd_sc_hd__decap_4 PHY_146 ();
 sky130_fd_sc_hd__decap_4 PHY_147 ();
 sky130_fd_sc_hd__decap_4 PHY_148 ();
 sky130_fd_sc_hd__decap_4 PHY_149 ();
 sky130_fd_sc_hd__decap_4 PHY_150 ();
 sky130_fd_sc_hd__decap_4 PHY_151 ();
 sky130_fd_sc_hd__decap_4 PHY_152 ();
 sky130_fd_sc_hd__decap_4 PHY_153 ();
 sky130_fd_sc_hd__decap_4 PHY_154 ();
 sky130_fd_sc_hd__decap_4 PHY_155 ();
 sky130_fd_sc_hd__decap_4 PHY_156 ();
 sky130_fd_sc_hd__decap_4 PHY_157 ();
 sky130_fd_sc_hd__decap_4 PHY_158 ();
 sky130_fd_sc_hd__decap_4 PHY_159 ();
 sky130_fd_sc_hd__decap_4 PHY_160 ();
 sky130_fd_sc_hd__decap_4 PHY_161 ();
 sky130_fd_sc_hd__decap_4 PHY_162 ();
 sky130_fd_sc_hd__decap_4 PHY_163 ();
 sky130_fd_sc_hd__decap_4 PHY_164 ();
 sky130_fd_sc_hd__decap_4 PHY_165 ();
 sky130_fd_sc_hd__decap_4 PHY_166 ();
 sky130_fd_sc_hd__decap_4 PHY_167 ();
 sky130_fd_sc_hd__decap_4 PHY_168 ();
 sky130_fd_sc_hd__decap_4 PHY_169 ();
 sky130_fd_sc_hd__decap_4 PHY_170 ();
 sky130_fd_sc_hd__decap_4 PHY_171 ();
 sky130_fd_sc_hd__decap_4 PHY_172 ();
 sky130_fd_sc_hd__decap_4 PHY_173 ();
 sky130_fd_sc_hd__decap_4 PHY_174 ();
 sky130_fd_sc_hd__decap_4 PHY_175 ();
 sky130_fd_sc_hd__decap_4 PHY_176 ();
 sky130_fd_sc_hd__decap_4 PHY_177 ();
 sky130_fd_sc_hd__decap_4 PHY_178 ();
 sky130_fd_sc_hd__decap_4 PHY_179 ();
 sky130_fd_sc_hd__decap_4 PHY_180 ();
 sky130_fd_sc_hd__decap_4 PHY_181 ();
 sky130_fd_sc_hd__decap_4 PHY_182 ();
 sky130_fd_sc_hd__decap_4 PHY_183 ();
 sky130_fd_sc_hd__decap_4 PHY_184 ();
 sky130_fd_sc_hd__decap_4 PHY_185 ();
 sky130_fd_sc_hd__decap_4 PHY_186 ();
 sky130_fd_sc_hd__decap_4 PHY_187 ();
 sky130_fd_sc_hd__decap_4 PHY_188 ();
 sky130_fd_sc_hd__decap_4 PHY_189 ();
 sky130_fd_sc_hd__decap_4 PHY_190 ();
 sky130_fd_sc_hd__decap_4 PHY_191 ();
 sky130_fd_sc_hd__decap_4 PHY_192 ();
 sky130_fd_sc_hd__decap_4 PHY_193 ();
 sky130_fd_sc_hd__decap_4 PHY_194 ();
 sky130_fd_sc_hd__decap_4 PHY_195 ();
 sky130_fd_sc_hd__decap_4 PHY_196 ();
 sky130_fd_sc_hd__decap_4 PHY_197 ();
 sky130_fd_sc_hd__decap_4 PHY_198 ();
 sky130_fd_sc_hd__decap_4 PHY_199 ();
 sky130_fd_sc_hd__decap_4 PHY_200 ();
 sky130_fd_sc_hd__decap_4 PHY_201 ();
 sky130_fd_sc_hd__decap_4 PHY_202 ();
 sky130_fd_sc_hd__decap_4 PHY_203 ();
 sky130_fd_sc_hd__decap_4 PHY_204 ();
 sky130_fd_sc_hd__decap_4 PHY_205 ();
 sky130_fd_sc_hd__decap_4 PHY_206 ();
 sky130_fd_sc_hd__decap_4 PHY_207 ();
 sky130_fd_sc_hd__decap_4 PHY_208 ();
 sky130_fd_sc_hd__decap_4 PHY_209 ();
 sky130_fd_sc_hd__decap_4 PHY_210 ();
 sky130_fd_sc_hd__decap_4 PHY_211 ();
 sky130_fd_sc_hd__decap_4 PHY_212 ();
 sky130_fd_sc_hd__decap_4 PHY_213 ();
 sky130_fd_sc_hd__decap_4 PHY_214 ();
 sky130_fd_sc_hd__decap_4 PHY_215 ();
 sky130_fd_sc_hd__decap_4 PHY_216 ();
 sky130_fd_sc_hd__decap_4 PHY_217 ();
 sky130_fd_sc_hd__decap_4 PHY_218 ();
 sky130_fd_sc_hd__decap_4 PHY_219 ();
 sky130_fd_sc_hd__decap_4 PHY_220 ();
 sky130_fd_sc_hd__decap_4 PHY_221 ();
 sky130_fd_sc_hd__decap_4 PHY_222 ();
 sky130_fd_sc_hd__decap_4 PHY_223 ();
 sky130_fd_sc_hd__decap_4 PHY_224 ();
 sky130_fd_sc_hd__decap_4 PHY_225 ();
 sky130_fd_sc_hd__decap_4 PHY_226 ();
 sky130_fd_sc_hd__decap_4 PHY_227 ();
 sky130_fd_sc_hd__decap_4 PHY_228 ();
 sky130_fd_sc_hd__decap_4 PHY_229 ();
 sky130_fd_sc_hd__decap_4 PHY_230 ();
 sky130_fd_sc_hd__decap_4 PHY_231 ();
 sky130_fd_sc_hd__decap_4 PHY_232 ();
 sky130_fd_sc_hd__decap_4 PHY_233 ();
 sky130_fd_sc_hd__decap_4 PHY_234 ();
 sky130_fd_sc_hd__decap_4 PHY_235 ();
 sky130_fd_sc_hd__decap_4 PHY_236 ();
 sky130_fd_sc_hd__decap_4 PHY_237 ();
 sky130_fd_sc_hd__decap_4 PHY_238 ();
 sky130_fd_sc_hd__decap_4 PHY_239 ();
 sky130_fd_sc_hd__decap_4 PHY_240 ();
 sky130_fd_sc_hd__decap_4 PHY_241 ();
 sky130_fd_sc_hd__decap_4 PHY_242 ();
 sky130_fd_sc_hd__decap_4 PHY_243 ();
 sky130_fd_sc_hd__decap_4 PHY_244 ();
 sky130_fd_sc_hd__decap_4 PHY_245 ();
 sky130_fd_sc_hd__decap_4 PHY_246 ();
 sky130_fd_sc_hd__decap_4 PHY_247 ();
 sky130_fd_sc_hd__decap_4 PHY_248 ();
 sky130_fd_sc_hd__decap_4 PHY_249 ();
 sky130_fd_sc_hd__decap_4 PHY_250 ();
 sky130_fd_sc_hd__decap_4 PHY_251 ();
 sky130_fd_sc_hd__decap_4 PHY_252 ();
 sky130_fd_sc_hd__decap_4 PHY_253 ();
 sky130_fd_sc_hd__decap_4 PHY_254 ();
 sky130_fd_sc_hd__decap_4 PHY_255 ();
 sky130_fd_sc_hd__decap_4 PHY_256 ();
 sky130_fd_sc_hd__decap_4 PHY_257 ();
 sky130_fd_sc_hd__decap_4 PHY_258 ();
 sky130_fd_sc_hd__decap_4 PHY_259 ();
 sky130_fd_sc_hd__decap_4 PHY_260 ();
 sky130_fd_sc_hd__decap_4 PHY_261 ();
 sky130_fd_sc_hd__decap_4 PHY_262 ();
 sky130_fd_sc_hd__decap_4 PHY_263 ();
 sky130_fd_sc_hd__decap_4 PHY_264 ();
 sky130_fd_sc_hd__decap_4 PHY_265 ();
 sky130_fd_sc_hd__decap_4 PHY_266 ();
 sky130_fd_sc_hd__decap_4 PHY_267 ();
 sky130_fd_sc_hd__decap_4 PHY_268 ();
 sky130_fd_sc_hd__decap_4 PHY_269 ();
 sky130_fd_sc_hd__decap_4 PHY_270 ();
 sky130_fd_sc_hd__decap_4 PHY_271 ();
 sky130_fd_sc_hd__decap_4 PHY_272 ();
 sky130_fd_sc_hd__decap_4 PHY_273 ();
 sky130_fd_sc_hd__decap_4 PHY_274 ();
 sky130_fd_sc_hd__decap_4 PHY_275 ();
 sky130_fd_sc_hd__decap_4 PHY_276 ();
 sky130_fd_sc_hd__decap_4 PHY_277 ();
 sky130_fd_sc_hd__decap_4 PHY_278 ();
 sky130_fd_sc_hd__decap_4 PHY_279 ();
 sky130_fd_sc_hd__decap_4 PHY_280 ();
 sky130_fd_sc_hd__decap_4 PHY_281 ();
 sky130_fd_sc_hd__decap_4 PHY_282 ();
 sky130_fd_sc_hd__decap_4 PHY_283 ();
 sky130_fd_sc_hd__decap_4 PHY_284 ();
 sky130_fd_sc_hd__decap_4 PHY_285 ();
 sky130_fd_sc_hd__decap_4 PHY_286 ();
 sky130_fd_sc_hd__decap_4 PHY_287 ();
 sky130_fd_sc_hd__decap_4 PHY_288 ();
 sky130_fd_sc_hd__decap_4 PHY_289 ();
 sky130_fd_sc_hd__decap_4 PHY_290 ();
 sky130_fd_sc_hd__decap_4 PHY_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_353 ();
endmodule
